���     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.3.0�ub�n_estimators�K�estimator_params�(hhhhhhhhhht��base_estimator��
deprecated��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h+�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Pclass��Sex��Age��SibSp��Parch��Fare��Embarked�et�b�n_features_in_�K�
n_outputs_�K�classes_�h*h-K ��h/��R�(KK��h4�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�
estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh&hNhJ�
hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h4�f8�����R�(KhMNNNJ����J����K t�b�C              �?�t�bhQh(�scalar���hLC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hK�
node_count�M�nodes�h*h-K ��h/��R�(KM��h4�V64�����R�(Kh8N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples��missing_go_to_left�t�}�(h}hLK ��h~hLK��hhLK��h�h]K��h�h]K ��h�hLK(��h�h]K0��h�h4�u1�����R�(Kh8NNNJ����J����K t�bK8��uK@KKt�b�B@E         �                     @"��p�?�           8�@    tati       u                    �?.y0��k�?�            �s@�d�X         "                    �?Hث3���?�            @m@ �P�X                             �?     ��?)             P@�P�X                          0�FF@�'N��?&            �N@       @                         s�,@�q�����?             9@      @������������������������       �                     @               	                 �܅3@8�A�0��?             6@        ������������������������       �                     @        
                        p�i@@�\��N��?             3@                                  �?��
ц��?	             *@                                   �?      �?             @        ������������������������       �                     �?                                  �H@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @                                  �<@և���X�?             @ �X  ������������������������       �                     @���X  ������������������������       �                     @P��X                             �?�q�q�?             @��X  ������������������������       �                     @P��X  ������������������������       �                      @���X                             �?�����H�?             B@��X  ������������������������       �                     9@���X                          p"�X@���|���?             &@��X                            �8@؇���X�?             @ ��X  ������������������������       �                     �?P��X  ������������������������       �                     @���X                             �?      �?             @ ��X  ������������������������       �                     �?���X  ������������������������       �                     @P��X          !                    �?�q�q�?             @��X  ������������������������       �                      @9F�X  ������������������������       �                     �?a��X  #       &                   �9@���Q��?i            @e@        $       %                    �?��s����?             5@        ������������������������       �                     @	X�X  ������������������������       �                     1@��X  '       f                  x#J@p�B<F]�?[            �b@
�X  (       G                     �?��c`��?L            �^@      0@)       >                   �>@8����?              G@)�X  *       +                    �?��
ц��?             :@ L�X  ������������������������       �                     @      @,       -                   �<@�q�q�?             5@ O�X  ������������������������       �                     @      �?.       =                    R@�<ݚ�?             2@�X  /       0                 03:@@�0�!��?             1@      @������������������������       �                     @MC�X  1       <                   �J@���!pc�?	             &@�X  2       3                 03k:@      �?              @ $�X  ������������������������       �                     �?      @4       ;                    H@����X�?             @��X  5       :                 X��B@r�q��?             @     �?6       7                 `fF<@      �?             @ �X  ������������������������       �                      @�G�X  8       9                 �|Y=@      �?              @ &�X  ������������������������       �                     �?�)�X  ������������������������       �                     �?�%�X  ������������������������       �                      @�M�X  ������������������������       �                     �?      @������������������������       �                     @       @������������������������       �                     �?��X  ?       @                 `f~I@ףp=
�?             4@&�X  ������������������������       �                     (@���X  A       B                 `��I@      �?              @ aram1 i������������������������       �                     �?      "CC       D                 03�I@؇���X�?             @    "eit������������������������       �                     �? name)
 E       F                    �?r�q��?             @ t_outpu������������������������       �                     �?or.
    ������������������������       �                     @ new_objH       e                    >@&:~�Q�?,             S@stimatoI       X                    �?�Y�R_�?+            �Q@ 

classJ       K                   @B@ �o_��?             9@  all es������������������������       �                     "@stimatorL       S                    -@     ��?             0@t the cM       P                   �'@      �?              @ argumenN       O                   �J@      �?              @ hod
   ������������������������       �                     �?es for t������������������������       �                     �?riginal Q       R                    D@�q�q�?             @        ������������������������       �                     @.__init_������������������������       �                      @explicitT       W                   �H@      �?              @ # intrU       V                   �E@      �?             @ ters
  ������������������������       �                      @gnature(������������������������       �                      @uding 's������������������������       �                     @r p in iY       d                    �?���}<S�?             G@= "selfZ       c                   @A@��-�=��?            �C@ paramet[       b                   �@@������?
             1@       \       ]                 �|Y=@�r����?	             .@ imators������������������������       �                     @meters i^       _                   �'@�<ݚ�?             "@(no var������������������������       �                     @sn't "
 `       a                 �|�=@�q�q�?             @ t_signa������������������������       �                      @ent name������������������������       �                     �?n parame������������������������       �                      @
       ������������������������       �                     6@        ������������������������       �                     @ If True������������������������       �                     @        g       t                 03�U@PN��T'�?             ;@s
     h       i                    <@��s����?             5@ mes map������������������������       �                     @      foj       k                    ?@      �?	             0@ attr(se������������������������       �                     �?ams") anl       m                    B@z�G�z�?             .@  = valu������������������������       �                     @ "__" + n       o                    C@�z�G��?             $@ value
 ������������������������       �                      @       "p       q                    �?      �?              @ od work������������������������       �                     @    (sucr       s                 0� Q@      �?             @ e
     ������������������������       �                     @o that i������������������������       �                     �?d object������������������������       �                     @s : dictv       w                    :@���B���?3            �S@    ----������������������������       �        
             1@tor instx                          �8@�jTM��?)            �N@ mple opy       ~                    @�g�y��?             ?@ turn sez       {                 ��W@      �?             @      ne������������������������       �                      @     for|       }                 �(\�?      �?              @ b_key =������������������������       �                     �?ams:
   ������������������������       �                     �?)
      ������������������������       �                     ;@d parame�       �                    �?��S���?             >@"Valid �       �                  DT@�ՙ/�?             5@       �       �                     �?�n_Y�K�?	             *@        �       �                 X�,D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�q�q�?             "@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 �UA@r�q��?             @       �       �                   @A@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 ���@�~�@
�?�            �x@        �       �                    7@�g�y��?             ?@        �       �                 03�@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     5@        �       
                ��Y7@�?��+�?�             w@       �       �                    /@����I�?�            �t@        �       �                    $@      �?             8@       ������������������������       �        	             .@        �       �                 �&�)@�q�q�?             "@        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        �       �                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?����Y��?�            s@        �       �                    �?���ȫ�?/            �T@        �       �                    �?�MI8d�?            �B@       �       �                    �?      �?             @@       ������������������������       �                     6@        �       �                  S�-@z�G�z�?             $@        ������������������������       �                      @        ������������������������       �                      @        �       �                 `�@1@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                     @X�<ݚ�?            �F@       �       �                  s@~�4_�g�?             F@        ������������������������       �                     @        �       �                   �3@      �?             D@        ������������������������       �                     �?        �       �                   �4@�99lMt�?            �C@        ������������������������       �                     @        �       �                 ��/@b�2�tk�?             B@       �       �                    �?�z�G��?             >@       �       �                   �5@�û��|�?             7@        ������������������������       �                     �?        �       �                    �?���|���?             6@       �       �                   P&@�q�q�?             5@       �       �                 �|�;@�z�G��?             4@       �       �                 pf�@�n_Y�K�?             *@        ������������������������       �                      @        �       �                 pf� @���!pc�?             &@       �       �                   �9@և���X�?             @       �       �                   �6@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ��� @؇���X�?             @       ������������������������       �                     @        �       �                  SE"@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?@�@+��?�            �k@        �       �                    �?�<ݚ�?             2@       �       �                   @@$�q-�?
             *@        �       �                 �|�:@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     "@        �       �                   �2@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�M��?}            �i@        �       �                    �?XB���?             =@       ������������������������       �                     <@        ������������������������       �                     �?        �       �                 �?�@h�V���?l             f@        �       �                   �?@�k~X��?.             R@       ������������������������       �        %             L@        �       �                   @@@      �?	             0@        �       �                   �@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                   �1@�ջ����?>             Z@        ������������������������       �                     (@        �       	                   �?��H�?7             W@       �                          �?z�G�z�?2            @U@       �       �                 @3�@*�s���?1             U@        �       �                   �?@      �?             ,@        �       �                   �9@�q�q�?             @       �       �                    �?      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �A@      �?              @        ������������������������       ��q�q�?             @        ������������������������       ����Q��?             @        �       �                   �2@؇���X�?*            �Q@        ������������������������       �                     @        �       �                 ��) @pH����?)            �P@        �       �                   �3@ 7���B�?             ;@        ������������������������       �                     �?        ������������������������       �                     :@        �       �                   �9@R���Q�?             D@        ������������������������       �                     1@        �                          (@��+7��?             7@       �                          ?@���Q��?             .@                              �|Y=@      �?              @        ������������������������       �                     @�aU�X                        �̜!@���Q��?             @ `U�X  ������������������������       �                     �?�_U�X                        �|�=@      �?             @ ^U�X  ������������������������       �                      @�]U�X  ������������������������       �                      @�\U�X  ������������������������       �                     @�[U�X  ������������������������       �                      @�ZU�X  ������������������������       �                     �?�YU�X  ������������������������       �                     @�XU�X                        ��T?@��-�=��?            �C@�zO�  ������������������������       �                     9@�zO�                           �?����X�?             ,@ �zO�  ������������������������       �                     @(�zO�                           @���|���?             &@�zO�                           @���Q��?             $@�zO�                        ��p@@�q�q�?             @ �zO�  ������������������������       �                     @�zO�  ������������������������       �                      @(�zO�  ������������������������       �                     @(�zO�  ������������������������       �                     �?(�zO�  �t�b�values�h*h-K ��h/��R�(KMKK��h]�BP        {@     Pq@     �`@      f@      ^@     �\@      2@      G@      1@      F@      *@      (@              @      *@      "@      @              $@      "@      @      @      @      @      �?               @      @              @       @              @      @              @      @              @       @      @                       @      @      @@              9@      @      @      �?      @      �?                      @      @      �?              �?      @              �?       @               @      �?             �Y@      Q@      1@      @              @      1@             @U@      P@     @T@     �D@      @@      ,@      ,@      (@              @      ,@      @              @      ,@      @      ,@      @      @               @      @      @      @              �?      @       @      @      �?      @      �?       @              �?      �?      �?                      �?       @                      �?      @                      �?      2@       @      (@              @       @              �?      @      �?      �?              @      �?              �?      @             �H@      ;@     �H@      6@      @      2@              "@      @      "@      @      @      �?      �?              �?      �?              @       @      @                       @       @      @       @       @               @       @                      @      E@      @     �A@      @      *@      @      *@       @      @              @       @      @              �?       @               @      �?                       @      6@              @                      @      @      7@      @      1@              @      @      (@      �?              @      (@              @      @      @       @              �?      @              @      �?      @              @      �?                      @      .@     �O@              1@      .@      G@      �?      >@      �?      @               @      �?      �?              �?      �?                      ;@      ,@      0@       @      *@       @      @      @      �?              �?      @              @      @              @      @                       @      @      @      �?       @      �?                       @      @      �?      @      �?              �?      @               @             �r@      Y@      >@      �?      "@      �?      "@                      �?      5@             �p@     �X@     @m@     �W@      @      5@              .@      @      @              @      @      �?       @              �?      �?      �?                      �?     �l@     �R@      ?@     �I@      @      ?@       @      >@              6@       @       @       @                       @      @      �?      @                      �?      9@      4@      9@      3@              @      9@      .@              �?      9@      ,@      @              6@      ,@      5@      "@      ,@      "@              �?      ,@       @      ,@      @      ,@      @       @      @               @       @      @      @      @      @      �?              �?      @                       @      @              @      �?      @              �?      �?              �?      �?                      �?              �?      @              �?      @      �?                      @              �?      i@      7@      ,@      @      (@      �?      @      �?       @              �?      �?      "@               @      @       @                      @     @g@      3@      <@      �?      <@                      �?     �c@      2@     �Q@      �?      L@              .@      �?      �?      �?              �?      �?              ,@             �U@      1@      (@             �R@      1@      Q@      1@     �P@      1@      @      @       @      @       @       @       @                       @               @      @      @       @      �?      @       @      N@      $@              @      N@      @      :@      �?              �?      :@              A@      @      1@              1@      @      "@      @       @      @              @       @      @              �?       @       @       @                       @      @               @              �?              @             �A@      @      9@              $@      @      @              @      @      @      @       @      @              @       @              @              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ/��hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtK�huh*h-K ��h/��R�(KK���h|�B�?                             @���*1�?�           8�@                                   @�7����?            �G@�R�X                              �?Pa�	�?            �@@ 5feb3c2                           �?z�G�z�?             @ 5.3"}@������������������������       �                     �?�aO�X  ������������������������       �                     @�bO�X  ������������������������       �                     <@�cO�X         	                 ��T?@؇���X�?             ,@ dO�X  ������������������������       �                      @        
                           @�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @               z                     @��?a�?�           ��@               !                    �?V$�݆��?�            �r@                                 0Cd=@Pns��ޭ?O            �`@                                  @E@$Q�q�?"            �O@                               ���*@p���?             I@                                `f�)@�IєX�?	             1@      ;@������������������������       �                     (@      "@                           :@z�G�z�?             @                                   5@      �?              @      @������������������������       �                     �?      @������������������������       �                     �?       @������������������������       �                     @       @������������������������       �                    �@@                                   �?�θ�?             *@     1@                        ���;@ףp=
�?             $@     (@������������������������       �                     "@      @������������������������       �                     �?                                   �?�q�q�?             @      G@������������������������       �                      @      �?������������������������       �                     �?      0@������������������������       �        -            �Q@        "       y                    �?4>���?t             e@      @#       8                 `ff:@�{��?��?n            @d@        $       '                    5@ >�֕�?0            �Q@      @%       &                   �2@      �?              @      �?������������������������       �                     �?      @������������������������       �                     �?        (       )                 �|Y=@ =[y��?.             Q@      @������������������������       �                     4@      �?*       7                   �*@      �?#             H@       +       ,                 `f�)@ȵHPS!�?             :@     @������������������������       �                     0@       @-       .                 �|�=@�z�G��?             $@      �?������������������������       �                     �?        /       4                   @D@�<ݚ�?             "@     �?0       3                   �A@؇���X�?             @        1       2                    @@�q�q�?             @       @������������������������       �                      @        ������������������������       �                     �?      @������������������������       �                     @        5       6                   �G@      �?              @      �?������������������������       �                     �?        ������������������������       �                     �?       @������������������������       �                     6@      �?9       V                    �?�)
;&��?>             W@        :       U                     �?�e����?            �C@     @;       T                   �H@��J�fj�?            �B@     �?<       Q                   @C@�g�y��?             ?@       =       >                   �4@�û��|�?             7@      "@������������������������       �                     @        ?       P                 �̾w@�G�z��?             4@      @@       M                    �?ҳ�wY;�?             1@     �?A       D                 �|�;@�q�q�?
             (@       @B       C                 Ȉ�P@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?      @E       L                   �A@�<ݚ�?             "@       F       K                 ��2>@�q�q�?             @        G       H                 `f&;@�q�q�?             @        ������������������������       �                     �?        I       J                 ���<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        N       O                   �7@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        R       S                 ���X@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        W       f                  i?@�c�����?"            �J@        X       e                   @>@p�ݯ��?             3@       Y       d                   �J@�t����?
             1@       Z       c                 `f�;@X�<ݚ�?             "@       [       ^                 �|�?@����X�?             @        \       ]                 �|�<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        _       `                   �C@z�G�z�?             @        ������������������������       �                     @        a       b                    H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        g       x                     �?@�0�!��?             A@       h       i                   �A@�n`���?             ?@        ������������������������       �                     "@        j       w                    �?���!pc�?             6@       k       v                    �?����X�?             5@       l       m                   �B@�z�G��?             4@        ������������������������       �                     @        n       u                 `f�K@@�0�!��?             1@       o       p                   �C@��S�ۿ?             .@       ������������������������       �                     "@        q       r                    �?r�q��?             @        ������������������������       �                     @        s       t                  x#J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        {       �                   �@@\�Yf�?�            �v@       |       �                    �?�8a�ME�?�            �s@        }       �                    �?@��Pl3�?<            @X@        ~       �                    �?     ��?             @@              �                    �?�>4և��?             <@       �       �                    �?�IєX�?             1@        ������������������������       �                      @        �       �                 �|�6@��S�ۿ?
             .@        ������������������������       �                     @        �       �                 ���@�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        �       �                    �?���|���?             &@        �       �                   �,@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?&����?(            @P@       �       �                 03�-@>���Rp�?%             M@       �       �                    �?�LQ�1	�?             G@       �       �                    �?8�Z$���?             :@       �       �                 ���@r�q��?             8@        ������������������������       �                     "@        �       �                   @@������?             .@       �       �                   �5@�q�q�?             "@        ������������������������       �                     �?        �       �                 �|=@      �?              @        ������������������������       �                      @        �       �                 �|�=@�q�q�?             @       ������������������������       �      �?             @        ������������������������       �                      @        �       �                 �|Y=@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 �|Y;@ףp=
�?             4@        ������������������������       �                     �?        �       �                  s�@�KM�]�?             3@        ������������������������       �                     @        �       �                    �?؇���X�?
             ,@       ������������������������       �8�Z$���?	             *@        ������������������������       �                     �?        �       �                 ��.@�q�q�?             (@        ������������������������       �                     @        �       �                 ��$1@և���X�?             @        ������������������������       �                     @        �       �                   �2@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�nYU}�?�             k@       �       �                    @�C�F��?o            �e@       �       �                 �|�=@�R����?n            �e@       �       �                    �?*~k���?b            �b@        �       �                  s@�eP*L��?             6@        ������������������������       �                     @        �       �                    4@�q�q�?             2@        �       �                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        �       �                 �|�;@d}h���?
             ,@       �       �                 pff@ףp=
�?             $@        �       �                   �7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                    �?x�]AgȽ?T             `@       �       �                    �?`Jj��?R             _@       �       �                 ���@�IєX�?N            �]@        �       �                   �5@����X�?             @        ������������������������       �                     @        �       �                 �&b@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                   �0@���>4ֵ?I             \@        �       �                 pFD!@      �?             @        ������������������������       �      �?              @        ������������������������       �                      @        �       �                 @3�!@ 7���B�?E             [@       �       �                 @3�@������?6            �T@       �       �                 �?$@���J��?!            �I@        �       �                 ��@���N8�?             5@       ������������������������       �        	             1@        �       �                 �|Y8@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @        ������������������������       �                     >@        �       �                 pf� @��a�n`�?             ?@       �       �                   �4@�8��8��?             8@        �       �                   �2@����X�?             @        ������������������������       �                      @        �       �                 0S5 @���Q��?             @       ������������������������       ��q�q�?             @        ������������������������       �                      @        ������������������������       �                     1@        �       �                    8@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     :@        �       �                 �Y�@z�G�z�?             @        ������������������������       �                      @        �       �                 pF�+@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   @@@8�A�0��?             6@       �       �                    �?      �?
             2@       �       �                    �?     ��?	             0@        ������������������������       �                     @        �       �                   �?@��
ц��?             *@        ������������������������       �                     @        �       �                 d�6@@���Q��?             $@       �       �                 ��I @և���X�?             @       �       �                 P�@      �?             @        ������������������������       �                      @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                 �̜2@d}h���?             E@        �       �                    <@�	j*D�?             *@       �       �                 P�@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     =@        ������������������������       �                     H@        �t�bh�h*h-K ��h/��R�(KK�KK��h]�B�       �{@     �p@      *@      A@      �?      @@      �?      @      �?                      @              <@      (@       @       @              @       @      @                       @     �z@     �m@     �a@     @d@      @      `@      @     �M@      �?     �H@      �?      0@              (@      �?      @      �?      �?              �?      �?                      @             �@@      @      $@      �?      "@              "@      �?               @      �?       @                      �?             �Q@      a@     �@@      `@     �@@     �P@      @      �?      �?      �?                      �?     @P@      @      4@             �F@      @      7@      @      0@              @      @              �?      @       @      @      �?       @      �?       @                      �?      @              �?      �?              �?      �?              6@             �O@      =@      7@      0@      5@      0@      .@      0@      ,@      "@      @              &@      "@      &@      @       @      @      �?       @               @      �?              @       @      @       @      �?       @              �?      �?      �?      �?                      �?      @              @              @       @               @      @                      @      �?      @              @      �?              @               @              D@      *@      (@      @      (@      @      @      @       @      @      �?      �?              �?      �?              �?      @              @      �?      �?      �?                      �?       @               @                       @      <@      @      9@      @      "@              0@      @      .@      @      ,@      @              @      ,@      @      ,@      �?      "@              @      �?      @              �?      �?      �?                      �?               @      �?              �?              @              @             �q@     �R@     �m@     �R@      N@     �B@      "@      7@      @      7@      �?      0@               @      �?      ,@              @      �?      &@      �?                      &@      @      @      @      �?              �?      @                      @      @             �I@      ,@      F@      ,@      D@      @      6@      @      4@      @      "@              &@      @      @      @              �?      @       @       @              @       @       @       @       @              @      �?              �?      @               @              2@       @      �?              1@       @      @              (@       @      &@       @      �?              @       @              @      @      @      @              �?      @      �?                      @      @             `f@      C@     @b@      =@     @b@      ;@     �`@      2@      (@      $@              @      (@      @      �?      @              @      �?              &@      @      "@      �?      �?      �?              �?      �?               @               @       @       @                       @     @^@       @      ]@       @      \@      @      @       @      @               @       @       @                       @     �Z@      @      @      �?      �?      �?       @              Z@      @     �S@      @      I@      �?      4@      �?      1@              @      �?      �?               @      �?      >@              <@      @      6@       @      @       @       @              @       @      �?       @       @              1@              @      �?      @                      �?      :@              @      �?       @               @      �?              �?       @              @              *@      "@      "@      "@      @      "@              @      @      @      @              @      @      @      @      �?      @               @      �?      �?      @                      @       @              @                       @     �@@      "@      @      "@       @      "@       @                      "@       @              =@              H@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJu�7hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�F         D                    �?���Yb�?�           8�@               )                    �?&ջ�{��?]            @b@      @                           �?JJ����?;            �W@       @                           �?��hJ,�?             A@    �M@������������������������       �                     ;@       @                        �ܙH@����X�?             @     9@������������������������       �                     @      @������������������������       �                      @       @	       
                   �2@      �?'             N@        ������������������������       �                     @                                     @����>4�?$             L@                                  @B@�ՙ/�?             5@                               ���<@      �?             0@        ������������������������       �                     @                                   �?�n_Y�K�?	             *@                               03SA@���Q��?             $@        ������������������������       �                     @                                @�6M@և���X�?             @      �?������������������������       �                     @                                X�,@@      �?             @                               �|Y<@      �?              @        ������������������������       �                     �?      @������������������������       �                     �?      �?������������������������       �                      @      @                        �nc@�q�q�?             @        ������������������������       �                     �?      @                        �̾w@      �?              @      @������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               "                 �|Y=@�#-���?            �A@     �R@        !                   @@z�G�z�?             $@     0@������������������������       �                      @        ������������������������       �                      @      >@#       $                 ���@`2U0*��?             9@ �X�X  ������������������������       �                     &@��X�X  %       (                 �|�=@@4և���?
             ,@�X�X  &       '                   @@      �?              @      @������������������������       �r�q��?             @0�X�X  ������������������������       �                      @0�X�X  ������������������������       �                     @0�X�X  *       3                     @R�}e�.�?"             J@�X�X  +       ,                    �?z�G�z�?             >@�X�X  ������������������������       �                     4@�X�X  -       2                    �?���Q��?             $@     �?.       1                     �?�q�q�?             @�X�X  /       0                 �U�X@z�G�z�?             @�X�X  ������������������������       �                     @��X�X  ������������������������       �                     �?      @������������������������       �                     �?p�X�X  ������������������������       �                     @      @4       =                    �?���|���?
             6@ �X�X  5       <                    �?և���X�?             ,@HX�X  6       9                    �?�eP*L��?             &@ �X�X  7       8                   �-@և���X�?             @ �X�X  ������������������������       �                     @��X�X  ������������������������       �                     @0�X�X  :       ;                 �|Y3@      �?             @ GX�X  ������������������������       �                     @��X�X  ������������������������       �                     �?0�X�X  ������������������������       �                     @��X�X  >       C                 03�-@      �?              @�X�X  ?       B                    �?�q�q�?             @     *@@       A                 �&�)@      �?              @ �X�X  ������������������������       �                     �?       @������������������������       �                     �?       ������������������������       �                     �?        ������������������������       �                     @      @E                       `f�S@��f
a�?r           ��@       F       �                 `f�$@�K�7���?]           Ȁ@        G       \                    �?��1��?�            �n@        H       S                   �6@�g�y��?             ?@        I       R                    �?r�q��?
             (@       J       O                    �?�<ݚ�?             "@       K       L                    �?؇���X�?             @        ������������������������       �                      @        M       N                   �3@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        P       Q                    4@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?       ������������������������       �                     @        T       Y                 ��@�d�����?             3@        U       V                 ���@�q�q�?             @        ������������������������       �                     �?        W       X                    �?z�G�z�?             @       ������������������������       �                     @       ������������������������       �                     �?       Z       [                    �?$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ]       b                   �0@d��]a��?�            �j@        ^       _                 pf�@���!pc�?             &@        ������������������������       �                     @        `       a                 pFD!@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        c       l                    �?����p�?�            �i@        d       e                 ���@�>4և��?             <@        ������������������������       �                      @        f       g                 �|Y=@      �?
             4@        ������������������������       �                     @       h       k                 X��A@�t����?	             1@       i       j                    �?؇���X�?             ,@       ������������������������       �8�Z$���?             *@       ������������������������       �                     �?       ������������������������       �                     @        m       �                 �|�=@����!p�?u             f@       n       {                 �?$@ ,V�ނ�?V            �_@        o       x                 ���@�L���?            �B@       p       q                     @�g�y��?             ?@        ������������������������       �                     "@        r       s                  Md@���7�?             6@        ������������������������       �                     &@        t       u                    7@�C��2(�?             &@        ������������������������       �                     @        v       w                   �8@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        y       z                 �|�;@�q�q�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @       |       �                    �?�x�E~�?;            @V@       }       �                    �?`���i��?:             V@       ~                        @3�@�D�e���?8            @U@        ������������������������       �                    �C@       �       �                   �;@�nkK�?             G@       �       �                   �9@�>����?             ;@       �       �                   �3@ ��WV�?             :@        �       �                   �2@�C��2(�?             &@        ������������������������       �                     @        �       �                 0S5 @؇���X�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �        	             .@        ������������������������       �                     �?        ������������������������       �                     3@        ������������������������       �                     @        ������������������������       �                     �?        �       �                   @@@ףp=
�?             I@        �       �                 �?�@�	j*D�?             *@        ������������������������       �                     @        �       �                    ?@X�<ݚ�?             "@        �       �                 �̌!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ��I @և���X�?             @       ������������������������       ����Q��?             @        ������������������������       �                      @        �       �                      @�?�|�?            �B@        ������������������������       �                     @        �       �                   �C@г�wY;�?             A@       �       �                   @C@�IєX�?             1@       ������������������������       �        
             .@        ������������������������       �      �?              @        ������������������������       �        	             1@        �       �                    �?��c���?�            0r@        �       �                    �?ڷv���?I            �\@        �       �                    �?Hm_!'1�?            �H@        ������������������������       �                     �?        �       �                    �?      �?             H@       �       �                     @ �Cc}�?             <@       �       �                     �?$�q-�?             :@        ������������������������       �                     @        �       �                   �A@�C��2(�?             6@       �       �                   �9@�IєX�?
             1@        �       �                   �'@؇���X�?             @        ������������������������       �                     @        �       �                   �3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        �       �                   �D@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ��&@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     4@        �       �                     @8�A�0��?*            �P@        �       �                     �?�}�+r��?             3@        ������������������������       �                     @        �       �                    �?��S�ۿ?             .@        �       �                    B@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             &@        �       �                    �?��k=.��?            �G@        ������������������������       �                      @        �       �                   @1@���V��?            �F@        �       �                    �?���|���?             &@       �       �                    D@����X�?             @       �       �                 �|�;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    0@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    @l��\��?             A@        �       �                    @����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    @ 7���B�?             ;@       ������������������������       �                     7@        �       �                   @D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �                          �?��|���?t             f@       �       �                    �?H%u��?T            @_@        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �       �                 `fF:@�S#א��?N            @]@       �       �                    4@����p�?+             Q@        �       �                    &@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        �       �                     @����˵�?$            �M@       �       �                   �*@���.�6�?             G@       �       �                 `f�)@ܷ��?��?             =@        ������������������������       �                     @        �       �                   �A@�LQ�1	�?             7@       �       �                    @@d}h���?             ,@       ������������������������       �                      @        ������������������������       �      �?             @        ������������������������       �                     "@        ������������������������       �                     1@        ������������������������       �                     *@        �                         �Q@Jm_!'1�?#            �H@       �                          �?r�q��?"             H@       �                             @t/*�?!            �G@       �       �                   �;@"pc�
�?             F@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �>@�p ��?            �D@        �       �                    K@     ��?             0@       �       �                   `G@�eP*L��?             &@       �       �                   @>@      �?              @       �       �                 `f�;@؇���X�?             @       �       �                 �|�<@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                  x#J@`2U0*��?             9@       ������������������������       �                     1@        �       �                 `�iJ@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?��[�8��?             �I@                                +@J�8���?             =@        ������������������������       �                     $@        ������������������������       �                     3@                                 @���7�?             6@       	      
                   �?      �?
             0@       ������������������������       �                     *@                                 @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                 �?�>4և��?             <@                                M@H%u��?             9@                              �k@�8��8��?             8@                               @E@�nkK�?             7@       ������������������������       �                     3@                                 �?      �?             @       ������������������������       �                     @       ������������������������       �                     �?        ������������������������       �                     �?       ������������������������       �                     �?                                 @�q�q�?             @        ������������������������       �                      @       ������������������������       �                     �?       �t�bh�h*h-K ��h/��R�(KMKK��h]�B�       �}@     �m@      P@     �T@      I@      F@      @      =@              ;@      @       @      @                       @     �F@      .@              @     �F@      &@      *@       @       @       @      @              @       @      @      @              @      @      @      @              �?      @      �?      �?              �?      �?                       @      �?       @              �?      �?      �?      �?                      �?      @              @@      @       @       @       @                       @      8@      �?      &@              *@      �?      @      �?      @      �?       @              @              ,@      C@      @      8@              4@      @      @       @      @      �?      @              @      �?              �?              @               @      ,@      @       @      @      @      @      @      @                      @      @      �?      @                      �?              @       @      @       @      �?      �?      �?              �?      �?              �?                      @     �y@     @c@     `y@     ``@     �j@     �@@      0@      .@       @      $@       @      @      �?      @               @      �?      @      �?                      @      �?      �?              �?      �?                      @      ,@      @       @      @      �?              �?      @              @      �?              (@      �?              �?      (@             �h@      2@       @      @      @              @      @              @      @             �g@      .@      7@      @       @              .@      @              @      .@       @      (@       @      &@       @      �?              @             �d@      $@     @^@      @      A@      @      >@      �?      "@              5@      �?      &@              $@      �?      @              @      �?              �?      @              @       @      @              �?       @     �U@       @     �U@       @     �T@       @     �C@              F@       @      9@       @      9@      �?      $@      �?      @              @      �?      �?      �?      @              .@                      �?      3@              @              �?             �F@      @      "@      @      @              @      @      �?      �?      �?                      �?      @      @       @      @       @              B@      �?      @             �@@      �?      0@      �?      .@              �?      �?      1@              h@     �X@     �E@      R@      @     �F@      �?              @     �F@      @      9@       @      8@              @       @      4@      �?      0@      �?      @              @      �?      �?      �?                      �?              $@      �?      @      �?                      @      �?      �?      �?                      �?              4@     �C@      ;@      �?      2@              @      �?      ,@      �?      @              @      �?                      &@      C@      "@               @      C@      @      @      @      @       @       @       @       @                       @      @               @       @               @       @              ?@      @      @       @      @                       @      :@      �?      7@              @      �?              �?      @             �b@      :@     �[@      .@      @      �?      @                      �?     �Y@      ,@     �O@      @      @       @               @      @              L@      @     �E@      @      :@      @      @              4@      @      &@      @       @              @      @      "@              1@              *@              D@      "@      D@       @     �C@       @      B@       @      �?       @              �?      �?      �?      �?                      �?     �A@      @      &@      @      @      @      @       @      @      �?      @      �?              �?      @              @                      �?              @      @              8@      �?      1@              @      �?              �?      @              @              �?                      �?      D@      &@      3@      $@              $@      3@              5@      �?      .@      �?      *@               @      �?       @                      �?      @              @      7@      @      6@       @      6@      �?      6@              3@      �?      @              @      �?              �?              �?               @      �?       @                      �?�t�bub�$>     hhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��!XhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM	huh*h-K ��h/��R�(KM	��h|�B@B         l                 ��%@�*���?�           8�@ �X                             /@,PY��?�             v@      "@������������������������       �                     @�'i�v,y5                        ���@j�q����?�            �u@ ���}��������������������������       �                    �E@    }t       3                 P�*@�A��t��?�            0s@  j           2                 �|Y>@J��D��?A             [@ j	           1                    �?���Q �?8            �X@     |	       
                 ��@r�qG�?7             X@        ������������������������       �                     �?                                  �?�|R���?6            �W@                                  �3@���B���?             :@                                �?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?�LQ�1	�?             7@                                  8@�C��2(�?             6@        ������������������������       �                     "@      ;@                        ��@8�Z$���?	             *@     "@                        ���@�C��2(�?             &@                                   �?�q�q�?             @      @������������������������       �                      @      @������������������������       �                     �?       @������������������������       �                      @       @                           @      �?              @        ������������������������       �                     �?     1@������������������������       �                     �?     (@������������������������       �                     �?      @       $                   �<@�㙢�c�?&            @Q@               #                   �6@�C��2(�?            �@@     G@                           �3@�S����?
             3@      �?������������������������       �                      @      0@!       "                    �?���!pc�?             &@        ������������������������       �                     @      @������������������������       �                      @        ������������������������       �                     ,@      @%       .                    �?      �?             B@     �?&       '                 ���@z�G�z�?             9@      @������������������������       �                      @        (       )                 �|Y=@�t����?             1@      @������������������������       �                     �?      �?*       +                 ���@      �?
             0@        ������������������������       ����Q��?             @     @,       -                 �Y�@�C��2(�?             &@       @������������������������       �                     @      �?������������������������       �      �?              @        /       0                 ��,@���|���?             &@     �?������������������������       �                     @        ������������������������       ��q�q�?             @       @������������������������       �                      @        ������������������������       �        	             $@      @4       i                    �?ȭ^���?x            �h@       5       <                 �?�@��ɉ�?v            `h@      �?6       ;                 �̌@�L#���?)            �P@        7       8                 �|Y=@���y4F�?             3@      @������������������������       �        
             *@      �?9       :                 ��]@�q�q�?             @        ������������������������       �                      @     @������������������������       �                     @     �?������������������������       �                     H@       =       B                     @     ��?M             `@      "@>       A                   �J@�+e�X�?             9@       ?       @                    �?�����?             3@       @������������������������       �                     @     �?������������������������       �                     *@�X�X  ������������������������       �                     @       @C       N                 @3�@�v�G���??            �Y@      @D       G                    �?      �?             0@ LX�X  E       F                   �9@���Q��?             @
Y�X  ������������������������       �                     @        ������������������������       �                      @p�X�X  H       I                    :@���|���?             &@        ������������������������       �                     @��X�X  J       K                   �?@և���X�?             @ Y�X  ������������������������       �                     �?p�X�X  L       M                   �A@      �?             @ �X�X  ������������������������       �      �?              @        ������������������������       �      �?             @pY�X  O       V                   �:@�=C|F�?4            �U@        P       U                   �3@`Ӹ����?            �F@ �X�X  Q       T                 0S5 @�����?
             5@ �X�X  R       S                   �1@�q�q�?             @ �X�X  ������������������������       �                     �?        ������������������������       �                      @��X�X  ������������������������       �                     2@��X�X  ������������������������       �                     8@p�X�X  W       X                   �;@d}h���?             E@        ������������������������       �                     @��X�X  Y       h                   �?@8�Z$���?            �C@       Z       [                 ��) @      �?             8@       ������������������������       �        	             &@        \       ]                   �<@��
ц��?             *@ �X�X  ������������������������       �                     @        ^       c                 P�*"@���Q��?             $@        _       `                 pf� @z�G�z�?             @ �X�X  ������������������������       �                      @��X�X  a       b                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        d       e                 ���"@���Q��?             @        ������������������������       �                      @        f       g                 �|Y=@�q�q�?             @  Y�X  ������������������������       �                      @        ������������������������       �                     �?0�X�X  ������������������������       �        	             .@pY�X  j       k                   �#@      �?             @ �X�X  ������������������������       �                      @�X�X  ������������������������       �                      @�X�X  m       �                  x#J@��d���?�            Pv@�X�X  n       �                    �?~���n��?�            Pp@        o       �                    @t�I��n�?R            @]@�X�X  p       u                    @f�����?N            �[@ HX�X  q       r                    @�}�+r��?             3@Y�X  ������������������������       �        
             0@        s       t                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @��X�X  v       �                     @ �&�T�?B             W@       w       �                   �H@�j��b�?(            �M@�X�X  x       �                    �?,�+�C�?%            �K@�X�X  y       z                     �?<���D�?            �@@ �X�X  ������������������������       �                     @0�X�X  {       �                   �7@8�Z$���?             :@�X�X  |       �                    �?������?             .@�X�X  }       �                    :@d}h���?             ,@ �X�X  ~                           �?      �?             @ Y�X  ������������������������       �                      @        ������������������������       �                      @0�X�X  �       �                    �?ףp=
�?	             $@        ������������������������       �                     �?        �       �                   �*@�����H�?             "@       �       �                 `f�)@؇���X�?             @        ������������������������       �                     �?        �       �                   �B@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     6@        �       �                 03�9@      �?             @       ������������������������       �                      @       ������������������������       �                      @        �       �                    �?4���C�?            �@@       �       �                 ��.@\X��t�?             7@       �       �                    �?�	j*D�?
             *@        �       �                 �|Y6@և���X�?             @       �       �                   �,@      �?             @        ������������������������       �                      @       �       �                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @       �       �                   �*@r�q��?             @        ������������������������       �                     �?       ������������������������       �                     @        �       �                    �?ףp=
�?             $@        ������������������������       �                     @        �       �                 �|Y>@r�q��?             @        ������������������������       �                     @        �       �                 03C3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 ���0@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@       ������������������������       �                     @       �       �                    @�q�q�?g             b@       �       �                    !@�θ�?^            @`@        ������������������������       �                     $@        �       �                 �&@r�q��?W             ^@        ������������������������       �                     �?       �       �                     �?�?��,�?V            �]@        �       �                 ��";@���j��?             G@        �       �                 ��$:@և���X�?
             ,@        ������������������������       �                     @        �       �                   �J@���!pc�?             &@       �       �                   @G@�����H�?             "@       �       �                    D@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     @       ������������������������       �                      @       �       �                    �?     ��?             @@       �       �                 ���=@�����?             5@        ������������������������       �                     $@       �       �                 p�i@@"pc�
�?             &@        �       �                 �|�;@�q�q�?             @        ������������������������       �                     �?        �       �                  �>@      �?              @        ������������������������       �                     �?       ������������������������       �                     �?       ������������������������       �                      @        �       �                   �<@���!pc�?	             &@        ������������������������       �                      @        �       �                 �|Y>@�����H�?             "@        �       �                 �|Y=@      �?             @        ������������������������       �                     �?       �       �                   �>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �*@�F��O�?8            @R@        �       �                   �@@�㙢�c�?             7@       ������������������������       �        
             (@        �       �                   �)@���|���?	             &@        ������������������������       �                      @        �       �                   �A@X�<ݚ�?             "@        ������������������������       �      �?             @        �       �                   @D@z�G�z�?             @        ������������������������       �                      @       �       �                    G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?`2U0*��?%             I@       �       �                 ��.@`Ql�R�?"            �G@        �       �                     @$�q-�?
             *@        ������������������������       �                     @        �       �                    �?r�q��?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     A@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             ,@        �                          @     ��?B             X@       �       �                    �?�n`���??            @W@       �       �                   �5@f>�cQ�?-            �N@        �       �                    �?X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @       �       �                    �?$�q-�?'             J@       �       �                      @�IєX�?&            �I@       �       �                   �B@ �q�q�?#             H@       �       �                    �?�IєX�?             A@       ������������������������       �                     <@        �       �                    �?�q�q�?             @       �       �                 X�,@@      �?             @       �       �                 p"�b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             ,@        �       �                 �|�;@�q�q�?             @        ������������������������       �                     �?        �       �                 �|�>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?       ������������������������       �                     �?                                �7@     ��?             @@                                 �?�C��2(�?             &@�zO�                           �?z�G�z�?             @ �zO�  ������������������������       �                     �?�zO�  ������������������������       �                     @(�zO�  ������������������������       �                     @�zO�                           �?�ՙ/�?             5@�zO�  ������������������������       �                     *@(�zO�  ������������������������       �                      @�zO�  ������������������������       �                     @(�zO�  �t�bh�h*h-K ��h/��R�(KM	KK��h]�B�       `|@     p@     �q@     �P@              @     �q@     �O@     �E@             �n@     �O@     �R@      A@      P@      A@      O@      A@              �?      O@     �@@      @      5@       @      �?              �?       @              @      4@       @      4@              "@       @      &@      �?      $@      �?       @               @      �?                       @      �?      �?      �?                      �?      �?             �L@      (@      >@      @      0@      @       @               @      @              @       @              ,@              ;@      "@      4@      @       @              (@      @              �?      (@      @       @      @      $@      �?      @              @      �?      @      @      @               @      @       @              $@             @e@      =@      e@      ;@     �O@      @      .@      @      *@               @      @       @                      @      H@             @Z@      7@      3@      @      *@      @              @      *@              @             �U@      1@      $@      @      @       @      @                       @      @      @      @              @      @              �?      @      @      �?      �?       @       @      S@      &@     �E@       @      3@       @      �?       @      �?                       @      2@              8@             �@@      "@              @     �@@      @      2@      @      &@              @      @      @              @      @      �?      @               @      �?       @               @      �?              @       @       @              �?       @               @      �?              .@               @       @               @       @             �d@     �g@     @b@     �\@      @@     @U@      :@     @U@      �?      2@              0@      �?       @      �?                       @      9@     �P@      @     �J@      @     �I@      @      =@              @      @      6@      @      &@      @      &@       @       @               @       @              �?      "@              �?      �?       @      �?      @              �?      �?      @              @      �?                       @      �?                      &@              6@       @       @               @       @              3@      ,@      $@      *@      "@      @      @      @      �?      @               @      �?      �?      �?                      �?      @              @      �?              �?      @              �?      "@              @      �?      @              @      �?      �?      �?                      �?      "@      �?              �?      "@              @             �\@      >@      Y@      >@              $@      Y@      4@              �?      Y@      3@     �@@      *@      @       @      @              @       @      �?       @      �?      @               @      �?       @              @       @              ;@      @      3@       @      $@              "@       @      �?       @              �?      �?      �?      �?                      �?       @               @      @               @       @      �?      @      �?      �?               @      �?              �?       @              @             �P@      @      3@      @      (@              @      @       @              @      @      �?      @      @      �?       @               @      �?              �?       @              H@       @      G@      �?      (@      �?      @              @      �?      @              �?      �?      �?                      �?      A@               @      �?              �?       @              ,@              5@     �R@      2@     �R@      "@      J@      @      @              @      @              @      H@      @      H@       @      G@       @      @@              <@       @      @      �?      @      �?      �?              �?      �?                       @      �?      �?              �?      �?                      ,@      �?       @              �?      �?      �?      �?                      �?      �?              "@      7@      �?      $@      �?      @      �?                      @              @       @      *@              *@       @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJC�NhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM	huh*h-K ��h/��R�(KM	��h|�B@B         p                     @���%&�?�           8�@    X         '                 �|Y=@N�ec�?�            ps@  l            
                 ��*@"��$�?G            �[@       @       	                    �?      �?             8@     �M@                           �?"pc�
�?             &@     @                        `f�)@�<ݚ�?             "@     E@������������������������       �                     @      @������������������������       �                      @      (@������������������������       �                      @      @������������������������       �        
             *@      @       "                 `fmj@�N��D�?6            �U@                                  �?���(\��?2             T@     �?                           6@�C��2(�?)            �P@                                   9@���|���?             &@       ������������������������       �                     @      0@                           �?z�G�z�?             @      @������������������������       �                     �?        ������������������������       �                     @      �?                           �?h㱪��?#            �K@       ������������������������       �                    �B@                                   �?�����H�?
             2@                                  5@��S�ۿ?             .@      @������������������������       �                     �?      �?������������������������       �                     ,@      @                           �?�q�q�?             @        ������������������������       �                     �?      @������������������������       �                      @      @                           �?d}h���?	             ,@                                   �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @     �R@        !                    �?���Q��?             @     0@������������������������       �                     @      @������������������������       �                      @        #       &                 0U�o@և���X�?             @     6@$       %                    5@z�G�z�?             @      ,@������������������������       �                     �?      @������������������������       �                     @      �?������������������������       �                      @        (       9                    �?4��@���?�             i@      @)       ,                    �?�nkK�?1            @Q@      �?*       +                 03�=@`2U0*��?             9@      >@������������������������       �                     �?      �?������������������������       �                     8@        -       6                    L@���7�?             F@      @.       /                   �B@��Y��]�?            �D@     @������������������������       �                     8@       @0       5                    -@�IєX�?             1@      �?1       2                   �'@�q�q�?             @      �?������������������������       �                     �?      �?3       4                    D@      �?              @      @������������������������       �                     �?      @������������������������       �                     �?      �?������������������������       �        	             ,@      �?7       8                   �L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        :       o                   �J@��ׂ�?Z            ``@     @;       n                 p�w@������?F            @Z@     H@<       a                   �G@��z6��?D             Y@     @=       >                   �)@� ���?6            @S@        ������������������������       �        	             ,@        ?       `                   �F@��s����?-            �O@     �?@       [                    �?�T`�[k�?(            �J@     7@A       L                    �?��Q���?             D@ �X�X  B       K                    �?     ��?
             0@      @C       J                    C@�q�q�?	             .@     @D       I                 ��2>@����X�?             ,@ LX�X  E       H                 ���<@      �?              @
Y�X  F       G                 ��";@z�G�z�?             @        ������������������������       �                     �?p�X�X  ������������������������       �                     @        ������������������������       �                     @��X�X  ������������������������       �                     @ Y�X  ������������������������       �                     �?p�X�X  ������������������������       �                     �? �X�X  M       Z                    �?      �?             8@       N       W                   @D@���!pc�?             6@Y�X  O       V                 `f�<@@�0�!��?             1@       P       U                 `fF:@���!pc�?             &@�X�X  Q       T                 `fv3@z�G�z�?             $@�X�X  R       S                 �|�=@����X�?             @ �X�X  ������������������������       �                      @        ������������������������       �                     @��X�X  ������������������������       �                     @��X�X  ������������������������       �                     �?p�X�X  ������������������������       �                     @        X       Y                     �?���Q��?             @ �X�X  ������������������������       �      �?              @       ������������������������       ��q�q�?             @       ������������������������       �                      @        \       ]                   �B@$�q-�?             *@ �X�X  ������������������������       �                     @        ^       _                 03�U@r�q��?             @       ������������������������       �                     @ �X�X  ������������������������       �                     �?��X�X  ������������������������       �                     $@        b       c                 `f4@
;&����?             7@        ������������������������       �                     @        d       i                    �?     ��?	             0@        e       f                    �?�q�q�?             @        ������������������������       �                      @  Y�X  g       h                 ���X@      �?             @       ������������������������       �                      @0�X�X  ������������������������       �                      @pY�X  j       k                 ���E@ףp=
�?             $@�X�X  ������������������������       �                      @�X�X  l       m                    �?      �?              @ �X�X  ������������������������       �                     �?�X�X  ������������������������       �                     �?        ������������������������       �                     @�X�X  ������������������������       �                     :@ HX�X  q                          @z6�>��?            y@Y�X  r       s                 ���@�o6�
�?�            �x@        ������������������������       �                     ;@        t                          @.�6�G,�?�             w@       u       �                    �?H?�߽��?�            �v@ �X�X  v       �                    �?�\��N��?H            �\@        w       |                    �?,���i�?            �D@�X�X  x       {                 ���@      �?             @@ �X�X  y       z                 0��@�q�q�?             @�X�X  ������������������������       �                      @0�X�X  ������������������������       �                     �?�X�X  ������������������������       �                     =@�X�X  }       ~                    @X�<ݚ�?             "@ �X�X  ������������������������       �                      @ Y�X         �                  S�2@և���X�?             @       �       �                    �?z�G�z�?             @ �X�X  ������������������������       �                      @        �       �                 ���&@�q�q�?             @        ������������������������       �                     �?       �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?       ������������������������       �                      @        �       �                    @:PZ(8?�?-            @R@        �       �                    @z�G�z�?             @        ������������������������       �                      @        �       �                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @       �       �                    ,@�t����?)             Q@        ������������������������       �                     $@        �       �                   �"@J�8���?$             M@        �       �                    @�ՙ/�?             5@       �       �                    ;@���Q��?             4@       �       �                    �?������?
             .@       �       �                 pf� @d}h���?	             ,@       �       �                   �7@�C��2(�?             &@        ������������������������       �                     @        �       �                 �&B@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @       �       �                    3@�q�q�?             @        ������������������������       �                     �?       ������������������������       �                      @        ������������������������       �                     �?        �       �                 �?� @z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 03�1@��G���?            �B@       �       �                    �?�X����?             6@       �       �                     @ҳ�wY;�?             1@       �       �                   �3@������?
             .@        ������������������������       �                     �?       �       �                   �0@d}h���?	             ,@       �       �                 �|�;@8�Z$���?             *@        ������������������������       �                      @        �       �                 ���.@���Q��?             @       �       �                    �?      �?             @       �       �                   �@@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?       ������������������������       �                      @       �       �                   �;@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@       �       �                 ��@H%u��?�            @o@        ������������������������       �                     @       �       �                    #@0�v����?�            �n@        �       �                     @     ��?             0@        ������������������������       �                     @        �       �                    @ףp=
�?             $@       �       �                    �?z�G�z�?             @        ������������������������       �                     �?        �       �                 ���A@      �?             @        �       �                    @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?,���>�?�            �l@        �       �                 03�-@д>��C�?'             M@       �       �                 �|Y=@ףp=
�?              I@        �       �                   �<@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        �       �                 �|Y?@��p\�?            �D@       �       �                    �?ܷ��?��?             =@       �       �                 ���@�����H�?             ;@        ������������������������       �                     @        �       �                 P�J@؇���X�?             5@       �       �                 ���@R���Q�?             4@        �       �                    �?�����H�?             "@       ������������������������       �r�q��?             @        ������������������������       �                     @       ������������������������       �"pc�
�?             &@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@       �       �                 ��.@      �?              @        ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                     �?       �       �                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �                         @@@���y�?p            �e@       �                          �?D��*�4�?\            @a@       �                          �?�[|x��?U            �_@       �       �                 �!&B@�H�@=��?M            �[@       �       �                 �|�=@ �h�7W�?J            �Z@       �       �                 @3�@��8�$>�?C            @X@       ������������������������       �        $             H@       �       �                 @�!@Hm_!'1�?            �H@       �       �                   � @PN��T'�?             ;@       �       �                 0S5 @�r����?             .@       �       �                   �3@؇���X�?             ,@        �       �                    1@�q�q�?             @        ������������������������       �                     �?       ������������������������       �                      @       ������������������������       �                     &@       ������������������������       �                     �?       �       �                   �7@r�q��?             (@       ������������������������       �                      @       �       �                 �|Y<@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     6@        �       �                   �?@�<ݚ�?             "@       �       �                   �>@���Q��?             @        �       �                 �̌!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 pff@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    ;@z�G�z�?             @        ������������������������       �                      @                                 >@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     .@        ������������������������       �                     (@        ������������������������       �                    �A@                               �:@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KM	KK��h]�B�       �{@     �p@     �`@      f@      <@     �T@      .@      "@       @      "@       @      @              @       @                       @      *@              *@     �R@      "@     �Q@      @      N@      @      @              @      @      �?              �?      @               @     �J@             �B@       @      0@      �?      ,@      �?                      ,@      �?       @      �?                       @      @      &@      �?       @      �?                       @       @      @              @       @              @      @      @      �?              �?      @                       @     �Z@     �W@      @     �P@      �?      8@      �?                      8@       @      E@      �?      D@              8@      �?      0@      �?       @              �?      �?      �?      �?                      �?              ,@      �?       @      �?                       @     �Y@      <@     @S@      <@     @S@      7@     @P@      (@      ,@             �I@      (@     �D@      (@      =@      &@      &@      @      $@      @      $@      @      @      @      @      �?              �?      @                      @      @                      �?      �?              2@      @      0@      @      ,@      @       @      @       @       @      @       @               @      @              @                      �?      @               @      @      �?      �?      �?       @       @              (@      �?      @              @      �?      @                      �?      $@              (@      &@      @              @      &@      @       @       @               @       @               @       @              �?      "@               @      �?      �?      �?                      �?              @      :@             0s@     @W@     �r@     @W@      ;@             0q@     @W@      q@     �V@      K@      N@      @      B@      �?      ?@      �?       @               @      �?                      =@      @      @               @      @      @      @      �?       @               @      �?      �?              �?      �?              �?      �?                       @     �H@      8@      �?      @               @      �?       @      �?                       @      H@      4@      $@              C@      4@       @      *@       @      (@      @      &@      @      &@      �?      $@              @      �?      @      �?                      @       @      �?              �?       @              �?              @      �?      @                      �?              �?      >@      @      .@      @      &@      @      &@      @              �?      &@      @      &@       @       @              @       @      @      �?      �?      �?              �?      �?               @                      �?              �?               @      @      �?              �?      @              .@             �k@      >@              @     �k@      ;@      "@      @              @      "@      �?      @      �?      �?              @      �?      �?      �?      �?                      �?       @              @             `j@      4@      H@      $@     �F@      @      @       @      @                       @      C@      @      :@      @      8@      @      @              2@      @      1@      @       @      �?      @      �?      @              "@       @      �?               @              (@              @      @              @      @       @              �?      @      �?      @                      �?     `d@      $@      `@      $@      ]@      $@     @Y@      $@      Y@      @     @W@      @      H@             �F@      @      7@      @      *@       @      (@       @      �?       @      �?                       @      &@              �?              $@       @       @               @       @               @       @              6@              @       @      @       @      �?      �?      �?                      �?       @      �?       @                      �?      @              �?      @               @      �?       @      �?                       @      .@              (@             �A@              �?      @              @      �?              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�R�[hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�C         \                    �?�s�ˈ.�?�           8�@               U                 p�H@�d�����?�            �l@ c a l        4                    �?Ҙ$�Ų�?k            �d@pñX                              @�<ݚ�?=            �X@  f e s        
                    �?�(\����?             D@  Param                          �J@�nkK�?             7@ handle������������������������       �                     4@
              	                 `f�2@�q�q�?             @ s
    -������������������������       �                     �?z�X  ������������������������       �                      @���X  ������������������������       �        
             1@VT�X                             �?:���W�?#            �M@ +�X                             �?�+e�X�?             9@ S�X                          H�%@���Q��?             $@ G�X  ������������������������       �                     @A{O�                          03�-@z�G�z�?             @ ��X  ������������������������       �                     @�"Y�X                          �|Y=@      �?              @      @������������������������       �                     �?        ������������������������       �                     �?p8Y�X                          X�,A@�r����?             .@+Y�X  ������������������������       �                     *@       @������������������������       �                      @      @       /                    �?�ʻ����?             A@     �?       .                    �?*;L]n�?             >@(Y�X                             '@П[;U��?             =@ :Y�X  ������������������������       �                     @      �?                          �4@      �?             :@ ;Y�X  ������������������������       �                     @      &@       )                 `��!@\X��t�?             7@      @       (                    C@������?	             .@      @        !                 P�@d}h���?             ,@ BY�X  ������������������������       �                     @      &@"       '                 �|Y>@      �?              @     �?#       &                 �|�;@      �?             @       $       %                   �8@      �?              @      @������������������������       �                     �?      @������������������������       �                     �?       @������������������������       �                      @      �?������������������������       �                     @        ������������������������       �                     �?       @*       +                    ;@      �?              @     @������������������������       �                     @      @,       -                   �@@�q�q�?             @      ;@������������������������       �                      @      @������������������������       �                     �?      @������������������������       �                     �?        0       1                    @      �?             @       @������������������������       �                     �?       @2       3                 ��l4@�q�q�?             @       @������������������������       �                     �?        ������������������������       �                      @      �?5       <                     @�'�=z��?.            �P@      �?6       9                    6@؇���X�?             5@       @7       8                 ��m1@      �?             @        ������������������������       �                      @      �?������������������������       �                      @      �?:       ;                   �B@�IєX�?             1@     "@������������������������       �                     0@      @������������������������       �                     �?      @=       @                    �?f.i��n�?            �F@      @>       ?                 ��.@�q�q�?             @      "@������������������������       �                      @      "@������������������������       �                     @        A       J                 03�1@��Sݭg�?            �C@ �X�X  B       I                    �?�q�q�?             (@      @C       H                 ��Y.@���Q��?             $@     @D       G                    �?z�G�z�?             @LX�X  E       F                    6@      �?             @ 
Y�X  ������������������������       �                     �?        ������������������������       �                     @p�X�X  ������������������������       �                     �?        ������������������������       �                     @��X�X  ������������������������       �                      @ Y�X  K       P                    @�>����?             ;@�X�X  L       O                 ���4@���7�?             6@ �X�X  M       N                 03C3@�q�q�?             @       ������������������������       �                      @Y�X  ������������������������       �                     �?       ������������������������       �        
             3@�X�X  Q       R                 ��T?@z�G�z�?             @ �X�X  ������������������������       �                      @ �X�X  S       T                    @�q�q�?             @        ������������������������       �                     �?��X�X  ������������������������       �                      @��X�X  V       [                 ���Q@$Q�q�?+            �O@ �X�X  W       X                    �?�J�4�?             9@       ������������������������       �                     3@ �X�X  Y       Z                 ���P@�q�q�?             @        ������������������������       �                      @       ������������������������       �                     @        ������������������������       �                     C@ �X�X  ]       �                    �?���A�
�?*           0~@        ^       k                 ��K.@N��c��?1            @S@        _       d                   �6@������?            �D@ �X�X  `       a                    �?      �?             @ �X�X  ������������������������       �                     �?        b       c                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        e       f                 �|=@�?�|�?            �B@        ������������������������       �                     &@  Y�X  g       j                   @@ ��WV�?             :@       h       i                 ���@�C��2(�?             &@�X�X  ������������������������       �                     @pY�X  ������������������������       �      �?             @�X�X  ������������������������       �                     .@�X�X  l       w                    �?b�2�tk�?             B@�X�X  m       r                 �|Y<@�z�G��?             4@ �X�X  n       q                    9@����X�?             @        o       p                    �?�q�q�?             @ �X�X  ������������������������       �                      @ HX�X  ������������������������       �                     �?Y�X  ������������������������       �                     @        s       v                   �F@$�q-�?
             *@        t       u                 X�,@@z�G�z�?             @       ������������������������       �                     @ �X�X  ������������������������       �                     �?        ������������������������       �                      @�X�X  x                           �?      �?             0@�X�X  y       |                 ��G@և���X�?
             ,@ �X�X  z       {                 ��3@      �?              @ �X�X  ������������������������       �                     @�X�X  ������������������������       �                     @�X�X  }       ~                 ���X@r�q��?             @�X�X  ������������������������       �                     @ Y�X  ������������������������       �                     �?       ������������������������       �                      @ �X�X  �       �                   �/@|g�&��?�            `y@,0,3,"K�       �                    �?<N_�U��?�            �p@�W�X  �       �                 �?�@     �?�             p@ �W�X  �       �                     @������?M            �^@ xW�X  ������������������������       �                     &@W",femal�       �                    �?�h����?E             \@ . Ander�       �                  ��@8�Z$���?             *@ 2,31.27������������������������       �                      @. 310130�       �                    �?"pc�
�?	             &@�W�X  �       �                 �|Y=@�<ݚ�?             "@ tW�X  ������������������������       �                     �?512,8.05�       �                 ��(@      �?              @|W�X  ������������������������       �r�q��?             @,,S
618,������������������������       �                      @male,26,������������������������       �                      @se",fema�       �                   �7@��:x�ٳ?:            �X@ e,26,0,������������������������       �                     A@��W�X  �       �                 �Yu@����?&            @P@1,0,117�       �                 �&B@(N:!���?            �A@653,15.�       �                   �8@`Jj��?             ?@ ,350029�       �                 �&b@���Q��?             @ TW�X  ������������������������       �                     @�:X�X  ������������������������       �                      @le,57,0,������������������������       �                     :@��W�X  �       �                    �?      �?             @ tcho",m������������������������       �                      @~W�X  ������������������������       �                      @on Henry������������������������       �                     >@��W�X  �       �                   �0@���H��?N            �`@ Maeglin�       �                 �̌!@�q�q�?             @ . Willi������������������������       �                      @�1X�X  ������������������������       �                     �?y",femal�       �                   �*@ ����?L            @`@",male,�       �                   �A@���5��?D            �\@8W�X  �       �                   �<@8�Z$���?7            �V@a (Mari�       �                   �3@$�q-�?             J@ ,"Thorn�       �                     @������?	             .@ Jensen,�       �                    &@      �?             @ �V�X  ������������������������       �      �?              @Skoog, M������������������������       �                      @,3,"Foo,�       �                   �1@���!pc�?             &@ Miss. E������������������������       �                     @`X�X  �       �                 0S5 @և���X�?             @ or, Mr.������������������������       �                     @ ?W�X  ������������������������       �                     @,3,"Will������������������������       �                    �B@P�W�X  �       �                 ��)"@��Sݭg�?            �C@X�X  �       �                   �?@�KM�]�?             3@Doling,�       �                   �>@8�Z$���?             *@ Mr. Jo�       �                 �|Y=@�8��8��?
             (@ _W�X  ������������������������       �                     �?�X�X  �       �                 ��) @�C��2(�?	             &@�U�X  ������������������������       �                     "@3.5,,S
6�       �                 pf� @      �?              @ �W�X  ������������������������       �                     �?5.5,,Q
6������������������������       �                     �?p8X�X  ������������������������       �                     �?.275,D48������������������������       �                     @�V�X  �       �                 �|�=@���Q��?             4@ �V�X  ������������������������       �                     @.5875,E5�       �                   �@@�t����?             1@�W�X  �       �                    $@�θ�?	             *@ �W�X  �       �                   �?@      �?             @ `W�X  ������������������������       �                     @P:W�X  ������������������������       �                     �?993,7.77������������������������       �                     "@,,S
670,������������������������       �      �?             @PpV�X  ������������������������       �                     7@�UW�X  ������������������������       �                     0@2,0,1,"D�       �                    �?���|���?             &@3,0,2,"�       �                     @X�<ݚ�?             "@ 7R�X  ������������������������       �                     �?`X�X  �       �                   �*@      �?              @ �W�X  �       �                 xFT$@���Q��?             @ 0,3,"Sa������������������������       �                      @ sW�X  ������������������������       �                     @
679,0,3������������������������       �                     @�W�X  ������������������������       �                      @PzW�X  �       �                    @4kMU*m�?X            `a@ �W�X  �       �                   �;@������?             .@ ,male,2������������������������       �                     @ Anderso�       �                    @      �?              @ s Edwar������������������������       �                     @s Willia������������������������       �                     @ nW�X  �                          �?���b��?P             _@:R�X  �       �                    �? �&�T�?:             W@<R�X  �       �                     @���3�E�?$             J@�V�X  �       �                 ��$:@�*/�8V�?             �G@ ,S
690,������������������������       �        	             .@�W�X  �       �                   �>@      �?             @@:W�X  �       �                 `fF<@�t����?             1@XW�X  �       �                    K@      �?             $@mW�X  �       �                 03k:@����X�?             @ �X  ������������������������       �                     �?��W�X  �       �                 �|�<@�q�q�?             @ ,male,4������������������������       �                      @�gW�X  �       �                 X��B@      �?             @ orland"������������������������       �                     �?P+X�X  �       �                   @G@�q�q�?             @1,1,"As������������������������       �      �?              @18,1,0,P������������������������       �                     �?ncer Vic������������������������       �                     @0�W�X  ������������������������       �                     @, Mr. Ma������������������������       �                     .@ iW�X  �       �                 �|�>@���Q��?             @ry Samu�       �                 �T�C@�q�q�?             @ 1,2,"Ke������������������������       �                     �?,,S
708,�       �                 �|�;@      �?              @ �W�X  ������������������������       �                     �?113781,1������������������������       �                     �?iam Geor������������������������       �                      @P�W�X  �       �                    �?      �?             D@�W�X  �       �                  x#J@r٣����?            �@@24,S
71������������������������       �        
             1@26,S
714�       �                    F@      �?             0@FX�X  �       �                 `f�K@�q�q�?             (@,0,3,"S�       �                    7@      �?              @ 8124,7.������������������������       �                     @��W�X  �       �                 `�iJ@z�G�z�?             @ ia ""Wi������������������������       �                      @��W�X  �       �                    @@�q�q�?             @ bW�X  ������������������������       �                      @Annie Je������������������������       �                     �?, Mr. Sv������������������������       �                     @�5X�X  ������������������������       �                     @, Mr. He�       �                 �|�:@����X�?             @ SW�X  ������������������������       �                     @vic, Mr.                            @�q�q�?             @  Peter ������������������������       �                     �?        ������������������������       �                      @                                 @      �?             @@                                �?`Jj��?             ?@                                 @�X�<ݺ?             2@        ������������������������       �                     @              
                   @@4և���?	             ,@             	                   0@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                 �?$�q-�?             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KMKK��h]�B�       �|@     @o@      N@      e@      L@     @[@      6@     @S@      �?     �C@      �?      6@              4@      �?       @      �?                       @              1@      5@      C@      @      3@      @      @              @      @      �?      @              �?      �?              �?      �?               @      *@              *@       @              .@      3@      *@      1@      *@      0@              @      *@      *@      @              $@      *@      @      &@      @      &@              @      @      @      @      �?      �?      �?      �?                      �?       @                      @      �?              @       @      @              �?       @               @      �?                      �?       @       @              �?       @      �?              �?       @              A@      @@      @      2@       @       @               @       @              �?      0@              0@      �?              ?@      ,@       @      @       @                      @      =@      $@      @       @      @      @      @      �?      @      �?              �?      @              �?                      @               @      9@       @      5@      �?       @      �?       @                      �?      3@              @      �?       @               @      �?              �?       @              @     �M@      @      5@              3@      @       @               @      @                      C@     y@     �T@     �M@      2@     �B@      @      �?      @              �?      �?       @               @      �?              B@      �?      &@              9@      �?      $@      �?      @              @      �?      .@              6@      ,@      ,@      @       @      @       @      �?       @                      �?              @      (@      �?      @      �?      @                      �?       @               @       @      @       @      @      @              @      @              �?      @              @      �?               @             `u@      P@      n@      :@     @m@      6@     @]@      @      &@             �Z@      @      &@       @       @              "@       @      @       @              �?      @      �?      @      �?       @               @             �W@      @      A@             �N@      @      ?@      @      =@       @      @       @      @                       @      :@               @       @               @       @              >@             @]@      0@      �?       @               @      �?              ]@      ,@      Y@      ,@     @S@      ,@      H@      @      &@      @      @      �?      �?      �?       @               @      @      @              @      @              @      @             �B@              =@      $@      1@       @      &@       @      &@      �?      �?              $@      �?      "@              �?      �?              �?      �?                      �?      @              (@       @              @      (@      @      $@      @      �?      @              @      �?              "@               @       @      7@              0@              @      @      @      @              �?      @      @       @      @       @                      @      @               @             @Y@      C@      @      &@              @      @      @              @      @             @X@      ;@     �P@      9@     �B@      .@     �A@      (@      .@              4@      (@      @      (@      @      @       @      @              �?       @      @               @       @       @      �?              �?       @      �?      �?              �?      @                      @      .@               @      @       @      �?      �?              �?      �?              �?      �?                       @      >@      $@      9@       @      1@               @       @      @       @      @      @      @              �?      @               @      �?       @               @      �?                      @      @              @       @      @              �?       @      �?                       @      >@       @      =@       @      1@      �?      @              *@      �?       @      �?              �?       @              @              (@      �?              �?      (@              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�v}hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtK�huh*h-K ��h/��R�(KK���h|�B@?         b                    �?��eC~�?�           8�@               ]                 p�H@������?�            `n@ u r n        D                    �?�H�]�r�?p            @e@     @       	                 ��@r�0p�?F            �Z@     @j@                           �?P���Q�?             4@       ������������������������       �        	             ,@                                ���@r�q��?             @     @������������������������       �                     @      �?������������������������       �                     �?      �?
                            @��V#�?8            �U@     �W@                           L@>A�F<�?             C@     8@                           �?     ��?             @@      0@������������������������       �                     @                                `f�)@�����H�?             ;@        ������������������������       �                     &@      7@                           �?     ��?             0@     (@                           :@r�q��?             (@ ��X  ������������������������       �                      @��X  ������������������������       �                     $@%�X                             <@      �?             @ |�X                            �9@      �?              @ ,�X  ������������������������       �                     �?�#�X  ������������������������       �                     �?<�X  ������������������������       �                      @��X                          `f�2@�q�q�?             @ �X  ������������������������       �                     @,��X  ������������������������       �                      @[	�X         7                 �|�<@     ��?              H@��X         ,                 Ь�!@�5��?             ;@#�X         #                   �6@���Q��?             .@ )�X         "                 �&B@�<ݚ�?             "@ �X          !                    4@      �?             @ ��X  ������������������������       �                      @      @������������������������       �                      @        ������������������������       �                     @     6@$       %                 �&B@�q�q�?             @      ,@������������������������       �                     �?      @&       '                   �9@���Q��?             @      �?������������������������       �                      @        (       )                   �@�q�q�?             @      @������������������������       �                     �?      �?*       +                 �?�@      �?              @      >@������������������������       �                     �?      �?������������������������       �                     �?        -       0                    �?r�q��?	             (@       @.       /                    4@�q�q�?             @      @������������������������       �                     �?       @������������������������       �                      @      �?1       6                 ��.@�����H�?             "@     �?2       3                   �-@z�G�z�?             @      �?������������������������       �                      @      @4       5                 �yG(@�q�q�?             @     @������������������������       �                      @      �?������������������������       �                     �?      �?������������������������       �                     @        8       =                 �|Y>@���N8�?             5@       9       :                    �?@4և���?             ,@       ������������������������       �                     $@     @;       <                    �?      �?             @      H@������������������������       �                     �?     @������������������������       �                     @        >       A                    @@և���X�?             @        ?       @                    �?      �?             @      �?������������������������       �                     �?     7@������������������������       �                     @       @B       C                   �A@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?      @E       J                    �?      �?*             P@        F       I                    �?���Q��?	             .@       G       H                 `�@1@�eP*L��?             &@        ������������������������       �                     @        ������������������������       �                     @       ������������������������       �                     @       K       L                    @Rg��J��?!            �H@        ������������������������       �                     @        M       N                    (@��6���?             E@        ������������������������       �                      @        O       P                   �:@�ʻ����?             A@        ������������������������       �        
             &@        Q       \                     @�LQ�1	�?             7@       R       [                    @X�<ݚ�?
             2@       S       T                   �?@��.k���?	             1@        ������������������������       �                     @        U       V                     @�q�q�?             (@        ������������������������       �                     @        W       X                    �?      �?              @        ������������������������       �                      @       Y       Z                 ��p@@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ^       _                    !@��pBI�?0            @R@        ������������������������       �                     �?        `       a                    @�k~X��?/             R@       ������������������������       �        .            �Q@        ������������������������       �                     �?        c       n                    @K�(i�?"           @}@        d       i                    �?8����?             7@       e       f                     @�q�q�?             (@       ������������������������       �                     @        g       h                 �y�-@����X�?             @        ������������������������       �                      @       ������������������������       �                     @       j       k                     @"pc�
�?             &@       ������������������������       �                     @       l       m                 pf�@@���Q��?             @        ������������������������       �                     @       ������������������������       �                      @        o       �                    �?4�<����?           �{@        p       {                 P�J.@����X�?4             U@        q       r                   @@     ��?             @@       ������������������������       �                     1@        s       z                 �(@z�G�z�?             .@        t       y                 �y�#@և���X�?             @       u       x                 �� @z�G�z�?             @       v       w                    ?@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @       |       �                    �?�E��
��?              J@       }       �                   �H@j���� �?            �I@       ~       �                     @      �?             E@              �                     �?��%��?            �B@       �       �                   �8@*;L]n�?             >@        �       �                  D�U@r�q��?             @ 01310,7������������������������       �                     �?.5,,Q
36������������������������       �                     @6,7.25,,�       �                    �?�q�q�?             8@n)",fem�       �                 �ܵ<@      �?             4@ oura Bo������������������������       �                      @ Annie",�       �                    �?r�q��?
             2@Pauline�       �                 `f�A@      �?             (@ George ������������������������       �                     @nd, Mr. �       �                 @�6M@      �?             @ an, Mr.������������������������       �                     @ghini, M������������������������       �                     @son, Mis������������������������       �                     @eyer, Mr�       �                 @��v@      �?             @8,,C
37������������������������       �                     @7077,7.2������������������������       �                     �?503,211.������������������������       �                     @.0125,,C�       �                    �?z�G�z�?             @ ,7.775,������������������������       �                     �?7,227.52������������������������       �                     @2,2653,1������������������������       �                     "@O 2. 310������������������������       �                     �?Mary Ali�       �                 `ff:@���5���?�            �v@ky, Mr.�       �                    �?��S�jC�?�            pr@harles �       �                    )@(�s���?�            �o@  Master������������������������       �                      @ss, Miss�       �                   @E@ ��GS=�?�            @o@atthew"�       �                   �D@�IєX�?�            �k@a",fema�       �                 ���@�X�<ݺ?�             k@ st",mal������������������������       �                    �C@ Olof",m�       �                 �?$@ ,��-�?i             f@ n Birge�       �                   �;@�㙢�c�?             7@ rjorie"������������������������       �                     @rs. Hjal�       �                    �?������?
             1@.7,G6,S�       �                 �|Y=@d}h���?             ,@ ,S
397,������������������������       �                      @
398,0,2������������������������       ��8��8��?             (@,2,"Pain�       �                 �|Y?@�q�q�?             @ Mrs. Wi������������������������       �                     �?3,"Niska������������������������       �                      @2,0,3,"A�       �                 �?�@�kb97�?[            @c@ la, Mis������������������������       �                    �A@rainen, �       �                   �3@T(y2��?C            �]@ 405,0,3�       �                   �1@��2(&�?             6@ 
406,0,������������������������       �                     @Widegren�       �                 0S5 @z�G�z�?	             .@ 1,2,"Ri�       �                   �2@      �?             @ 09,0,3,������������������������       �                     �?.775,,S
������������������������       ��q�q�?             @
411,0,3������������������������       �                     &@,"Hart, �       �                    �?h�a��?7            @X@iss. Da�       �                 �|�=@ rpa�?5            @W@Mr. Alf�       �                 @3�!@��v$���?!            �N@ Johan J�       �                 pf� @�nkK�?             7@ek, Mrs������������������������       �        
             4@,S
417,1�       �                    8@�q�q�?             @ le,34,1������������������������       �                      @,female,������������������������       �                     �?,male,30������������������������       �                     C@ale,10,0�       �                   �?@      �?             @@ ,0,0,34�       �                     @�<ݚ�?             "@ A/5. 13������������������������       �                     @15082,7.�       �                 @3�@      �?             @ aria Br������������������������       �                     �?r. Vikto�       �                 �̌!@�q�q�?             @ , Mr. P������������������������       �                      @Mrs. Cha������������������������       �                     �?8,1,2,"P�       �                   �@@���}<S�?             7@ Marshal������������������������       �                     "@es",male�       �                     @؇���X�?	             ,@mbisky)�       �                   �3@؇���X�?             @strom-S�       �                   �A@r�q��?             @ 52,S
43������������������������       ��q�q�?             @",female������������������������       �                     @der (Ali������������������������       �                     �?3,"Kalli�       �                 @3�@؇���X�?             @ 5,,S
43������������������������       ��q�q�?             @,E44,S
4������������������������       �                     @120,B96 ������������������������       �                     @emale,21�       �                 ���%@z�G�z�?             @ (Emily ������������������������       �                     @ Mr. Mar������������������������       �      �?              @, Mr. Jo������������������������       �                     =@41,1,2,"�       �                     @ qP��B�?            �E@ 1,F.C.C������������������������       �                      @45769,9.�       �                   �/@��?^�k�?            �A@76,7.77������������������������       �                     2@30434,13�       �                    )@�IєX�?             1@ ,65306,������������������������       �                     �?,33638,8������������������������       �        
             0@,female,�       �                    �?:ɨ��?-            �P@r",male�       �                    �?���Q��?              I@herine"�       �                     �?��.k���?             A@thur Go�       �                   �>@X�<ݚ�?             ;@Edwy Ar�       �                    R@����X�?             5@r. Ingv�       �                   @=@�q�q�?             2@an, Mr.�       �                 �|�<@���Q��?             $@ 1,1,"Go������������������������       �                     �?455,0,3,�       �                 `f�;@�q�q�?             "@"Jalsev�       �                 �|�?@      �?              @ t, Mr. ������������������������       �                     @nyon, Mr�       �                   �J@���Q��?             @ 459,1,2������������������������       �                     @S
460,0,������������������������       �                      @,1,"Ande������������������������       �                     �?Morley, ������������������������       �                      @. Arthur������������������������       �                     @Jacob Ch������������������������       �                     @Simon",m�       �                 �|�>@؇���X�?             @Estansl������������������������       �                     @bell, Mr������������������������       �                     �?n Montgo�       �                 ��9L@      �?
             0@ames",m�       �                   �C@ףp=
�?             $@ rbara",������������������������       �                     @ur",male�       �                    G@�q�q�?             @0,31508�       �                     �?      �?              @ th)",fe������������������������       �                     �?in S (Ma������������������������       �                     �?7917,D,C������������������������       �                     �?3,9.8375�       �                   �D@      �?             @5,52,A1�       �                     �?      �?             @1,,S
47������������������������       �                     @8,,S
479������������������������       �                     �?08,,S
48������������������������       �                      @.2875,,S������������������������       �                     0@2144,46.�t�b��     h�h*h-K ��h/��R�(KK�KK��h]�B�       p|@      p@     �O@     �f@     �N@     @[@      =@     @S@      �?      3@              ,@      �?      @              @      �?              <@      M@      @      ?@      @      =@              @      @      8@              &@      @      *@       @      $@       @                      $@      �?      @      �?      �?              �?      �?                       @      @       @      @                       @      5@      ;@      0@      &@      @      "@       @      @       @       @       @                       @              @      @       @      �?              @       @       @              �?       @              �?      �?      �?      �?                      �?      $@       @       @      �?              �?       @               @      �?      @      �?       @               @      �?       @                      �?      @              @      0@      �?      *@              $@      �?      @      �?                      @      @      @      @      �?              �?      @              �?       @               @      �?              @@      @@      "@      @      @      @      @                      @      @              7@      :@              @      7@      3@       @              .@      3@              &@      .@       @      $@       @      "@       @      @              @       @              @      @      @       @               @      @              @       @              �?              @               @     �Q@      �?              �?     �Q@             �Q@      �?             �x@      S@      @      0@      @      @              @      @       @               @      @               @      "@              @       @      @              @       @             x@      N@      N@      8@      =@      @      1@              (@      @      @      @      @      �?       @      �?              �?       @               @                       @       @              ?@      5@      >@      5@      5@      5@      4@      1@      *@      1@      @      �?              �?      @               @      0@      @      .@       @              @      .@      @      "@              @      @      @      @                      @              @      @      �?      @                      �?      @              �?      @      �?                      @      "@              �?             Pt@      B@     pq@      0@     �m@      .@               @     �m@      *@      j@      *@     �i@      (@     �C@             �d@      (@      3@      @      @              *@      @      &@      @               @      &@      �?       @      �?              �?       @             @b@       @     �A@             �[@       @      3@      @      @              (@      @      �?      @              �?      �?       @      &@              W@      @      V@      @      N@      �?      6@      �?      4@               @      �?       @                      �?      C@              <@      @      @       @      @               @       @              �?       @      �?       @                      �?      5@       @      "@              (@       @      @      �?      @      �?       @      �?      @              �?              @      �?       @      �?      @              @              @      �?      @              �?      �?      =@              E@      �?       @              A@      �?      2@              0@      �?              �?      0@              G@      4@      >@      4@      2@      0@      (@      .@      @      .@      @      (@      @      @              �?      @      @      @      @      @               @      @              @       @              �?                       @              @      @              @      �?      @                      �?      (@      @      "@      �?      @               @      �?      �?      �?              �?      �?              �?              @      @      �?      @              @      �?               @              0@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJg}�XhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMChuh*h-K ��h/��R�(KMC��h|�B�P         r                 `f�$@��t���?�           8�@                                    @z�G�z�?�            @p@       @������������������������       �                      @�'i�v,y5       k                   @@@Z���c��?�            �o@���}��                            �?�۲I <�?�            �j@      @                        �|Y=@T�7�s��?#            �L@       @                        ���@"pc�
�?             &@      ;@       	                   �2@�q�q�?             @       @������������������������       �                     �?        
                        �{@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                03@�LQ�1	�?             G@                               ���@���"͏�?            �B@                                   �?$�q-�?             *@        ������������������������       �                     �?      �?������������������������       �                     (@                                   �?�q�q�?             8@     �?                        ��@�LQ�1	�?             7@        ������������������������       �                      @      �?                           �?����X�?             5@     3@                           �?�q�q�?             2@      C@������������������������       �                     @      @                        ���@؇���X�?	             ,@        ������������������������       �                     �?      �?������������������������       �8�Z$���?             *@      ,@������������������������       �                     @        ������������������������       �                     �?      �?                           �?�<ݚ�?             "@      @������������������������       �                     @        ������������������������       �                      @        !       4                    �?�IA��?e            �c@      0@"       3                 �|Y>@     ��?             0@     "@#       2                    �?���Q��?             .@     @$       -                   �6@և���X�?             ,@     �?%       ,                 xF� @X�<ݚ�?             "@     @&       +                    �?r�q��?             @     0@'       *                   �3@z�G�z�?             @      *@(       )                 P��@      �?              @      @������������������������       �                     �?       @������������������������       �                     �?        ������������������������       �                     @      @������������������������       �                     �?      �?������������������������       �                     @      @.       /                 �&B@z�G�z�?             @      �?������������������������       �                      @      @0       1                    9@�q�q�?             @     �?������������������������       �                      @       @������������������������       �                     �?      �?������������������������       �                     �?      �?������������������������       �                     �?      �?5       H                 �?�@`	�<��?V            �a@     �?6       E                   �?@��p\�?.            �T@     �?7       <                 ���@ �\���?,            �S@      4@8       9                    7@����X�?             @      (@������������������������       �                     @      @:       ;                 �&b@      �?             @       ������������������������       �                      @        ������������������������       �                      @      @=       D                 �?$@������?'             R@      �?>       ?                 �|Y;@HP�s��?             9@     @������������������������       �        
             2@        @       C                 �|Y>@����X�?             @       A       B                 ��@���Q��?             @      @������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @      @������������������������       �                    �G@        F       G                   �@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        I       R                 @3�@��$�4��?(            �M@        J       Q                    �?X�<ݚ�?             "@       K       P                    �?      �?              @       L       M                   �9@և���X�?             @        ������������������������       �                      @        N       O                   �?@���Q��?             @        ������������������������       �                     �?        ������������������������       �      �?             @        ������������������������       �                     �?       ������������������������       �                     �?       S       h                 �|�=@j�q����?"             I@       T       a                 @�!@��0{9�?             �G@       U       ^                   � @"pc�
�?            �@@       V       ]                 0S5 @�>4և��?             <@       W       \                   �4@�+$�jP�?             ;@        X       Y                    1@X�<ݚ�?             "@        ������������������������       �      �?             @        Z       [                   �2@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @        ������������������������       �                     2@        ������������������������       �                     �?        _       `                   �7@z�G�z�?             @       ������������������������       �                     @       ������������������������       �                     �?        b       c                 ���"@@4և���?
             ,@        ������������������������       �                     @        d       e                   �<@ףp=
�?             $@       ������������������������       �                     @       f       g                 �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @       i       j                    ?@�q�q�?             @        ������������������������       �                      @       ������������������������       �                     �?       l       m                   @C@P�Lt�<�?             C@        ������������������������       �                     3@       n       o                    �?�}�+r��?             3@        ������������������������       �                      @        p       q                   �C@�IєX�?
             1@        ������������������������       ��q�q�?             @       ������������������������       �                     ,@        s                           @.iI\��?           0|@       t       �                  x#J@$;hB��?�            @s@       u       �                   �<@��U��?�            �j@        v       �                    �?��V#�?1            �U@       w       x                    �?@3����?             K@        ������������������������       �                      @        y       �                    �?��<b�ƥ?             G@        z       {                   �6@�nkK�?	             7@        ������������������������       �                     "@       |                          �9@@4և���?             ,@        }       ~                    �?z�G�z�?             @        ������������������������       �                     �?       ������������������������       �                     @       ������������������������       �                     "@        ������������������������       �                     7@ 01310,7�       �                    �?     ��?             @@ 5,,Q
36�       �                    �?և���X�?             @,7.25,,�       �                   �8@���Q��?             @n)",fem�       �                 hf:@�q�q�?             @ oura Bo������������������������       �                      @ Annie",������������������������       �                     �?Pauline������������������������       �                      @ George ������������������������       �                      @nd, Mr. �       �                   �>@HP�s��?             9@an, Mr.������������������������       �                     7@ghini, M������������������������       �                      @son, Mis�       �                    �?b����?R            �_@yer, Mr�       �                  �?@�8�Վ��?Q            @_@8,,C
37�       �                    �?D��ٝ�?B            @Y@ 077,7.2�       �                    �?�eP*L��?             6@ 03,211.�       �                    D@r�q��?             @0125,,C������������������������       �                     @ ,7.775,������������������������       �                     �?7,227.52�       �                   @C@     ��?	             0@,2653,1�       �                 ��";@r�q��?             (@ 2. 310�       �                   @@@�q�q�?             @ ary Ali������������������������       �                     @ky, Mr.�       �                   �A@�q�q�?             @ harles ������������������������       �                      @  Master������������������������       �                     �?ss, Miss������������������������       �                     @atthew"�       �                     �?      �?             @ a",fema������������������������       �                     @ st",mal������������������������       �                     �? Olof",m�       �                    �?���%&�?5            �S@n Birge�       �                   �F@^H���+�?2            �R@rjorie"�       �                   @F@�[�IJ�?             �G@s. Hjal�       �                   @E@�lg����?            �E@.7,G6,S�       �                     �?�e����?            �C@ ,S
397,�       �                 �|�?@�q�q�?             @398,0,2�       �                   �>@z�G�z�?             @2,"Pain�       �                 `f�;@      �?              @ Mrs. Wi������������������������       �                     �?3,"Niska������������������������       �                     �?2,0,3,"A������������������������       �                     @ la, Mis������������������������       �                     �?rainen, �       �                   �C@4���C�?            �@@405,0,3�       �                   @B@����"�?             =@
406,0,�       �                    �?
;&����?             7@ idegren������������������������       �                     "@ 1,2,"Ri�       �                    1@؇���X�?             ,@09,0,3,�       �                   �'@�<ݚ�?             "@ 775,,S
������������������������       �                     @
411,0,3�       �                    @@�q�q�?             @ "Hart, ������������������������       �                     @iss. Da������������������������       ��q�q�?             @Mr. Alf������������������������       �                     @ Johan J������������������������       �                     @ek, Mrs�       �                   �,@      �?             @ S
417,1������������������������       �      �?              @ le,34,1������������������������       �                      @,female,������������������������       �                     @,male,30������������������������       �                     @ale,10,0�       �                   �R@�<ݚ�?             ;@,0,0,34�       �                    �?���B���?             :@ A/5. 13������������������������       �                     @15082,7.�       �                    �?���}<S�?             7@aria Br�       �                   �I@�C��2(�?             6@. Vikto�       �                 ��:@r�q��?             (@, Mr. P������������������������       �                      @Mrs. Cha�       �                 `f�;@      �?             @,1,2,"P������������������������       �                      @ Marshal������������������������       �                      @es",male������������������������       �                     $@mbisky)������������������������       �                     �?strom-S������������������������       �                     �? 52,S
43�       �                    �?z�G�z�?             @ ,female������������������������       �                     �?der (Ali������������������������       �                     @3,"Kalli�       �                    �?      �?             8@ 5,,S
43������������������������       �                     @,E44,S
4������������������������       �                     5@120,B96 ������������������������       �                     �?emale,21�                         �O@�q�q�?A             X@(Emily �       �                   �5@���!pc�?>             V@ Mr. Mar�       �                   �1@��.k���?             1@ Mr. Jo�       �                 ��f`@؇���X�?             @1,1,2,"������������������������       �                     @ 1,F.C.C�       �                    �?      �?              @ 5769,9.������������������������       �                     �?76,7.77������������������������       �                     �?30434,13�       �                    �?z�G�z�?             $@,65306,������������������������       �                      @,33638,8������������������������       �                      @,female,�       �                 `fmj@@���?T�?3            �Q@r",male�       �                    �?     8�?.             P@herine"�       �                 ���P@���-T��?-             O@ thur Go�       �                 03sP@�z�G��?             4@Edwy Ar�       �                    �?@�0�!��?             1@ r. Ingv������������������������       �                     $@an, Mr.�       �                   �H@և���X�?             @1,1,"Go�       �                    �?z�G�z�?             @ 55,0,3,������������������������       �                     @"Jalsev�       �                 0�nL@      �?              @ t, Mr. ������������������������       �                     �?nyon, Mr������������������������       �                     �? 459,1,2������������������������       �                      @S
460,0,������������������������       �                     @,1,"Ande�       �                    �?@4և���?              E@orley, �       �                    �?@-�_ .�?            �B@ Arthur�       �                    �?`Jj��?             ?@acob Ch������������������������       �                     0@Simon",m�       �                    �?�r����?             .@ Estansl������������������������       �                     @bell, Mr�       �                   �H@      �?              @ Montgo�       �                 ЈT@؇���X�?             @ ames",m������������������������       �                     @ rbara",�       �                   �D@      �?             @ r",male������������������������       �                      @0,31508�       �                 Ј�U@      �?              @ th)",fe������������������������       �                     �?in S (Ma������������������������       �                     �?7917,D,C������������������������       �                     �?3,9.8375������������������������       �                     @5,52,A1�       �                 ��W@z�G�z�?             @ 1,,S
47������������������������       �                     @8,,S
479������������������������       �                     �?08,,S
48������������������������       �                      @.2875,,S�       �                    �?և���X�?             @ 144,46.������������������������       �                     �?0,0,2398�                          �?      �?             @5 3594,                       �̾w@���Q��?             @34,9.58������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @                                 �?x�f��^�?[            �a@                                 �?�>$�*��?            �D@                             X�,A@��+7��?             7@             	                  �0@��s����?             5@        ������������������������       �                     @        
                        �7@������?             .@        ������������������������       �                     �?                              �|Y=@d}h���?             ,@        ������������������������       �                      @                                 �?      �?             (@                              S�-@�z�G��?             $@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @                                 �?�q�q�?             2@                             03�-@�eP*L��?             &@                                 3@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                 �?r�q��?             @                                �2@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @              8                   �?t�F�}�?B            �Y@              /                   �?�q�q�?'             N@        !      *                ���5@*;L]n�?             >@       "      )                  �D@     ��?
             0@       #      (                   7@�r����?	             .@        $      '                   �?      �?             @       %      &                   +@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        +      .                  @C@����X�?             ,@        ,      -                X��@@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        0      1                   )@������?             >@        ������������������������       �                     @        2      7                   ;@H%u��?             9@        3      6                   �?և���X�?             @        4      5                �!&B@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     2@        9      B                   @@4և���?             E@        :      ;                   �?���!pc�?             &@        ������������������������       �                     @        <      =                   @և���X�?             @        ������������������������       �                     @        >      ?                   �?      �?             @        ������������������������       �                      @        @      A                ��T?@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ?@        �t�bh�h*h-K ��h/��R�(KMCKK��h]�B0       �{@     �p@      j@      J@       @              i@      J@     `d@     �I@      @@      9@       @      "@       @      �?      �?              �?      �?      �?                      �?               @      >@      0@      <@      "@      (@      �?              �?      (@              0@       @      .@       @               @      .@      @      (@      @              @      (@       @      �?              &@       @      @              �?               @      @              @       @             ``@      :@      "@      @      "@      @       @      @      @      @      �?      @      �?      @      �?      �?              �?      �?                      @              �?      @              @      �?       @               @      �?       @                      �?      �?                      �?     �^@      3@      S@      @     �R@      @      @       @      @               @       @       @                       @     �Q@       @      7@       @      2@              @       @      @       @      @                       @       @             �G@              �?       @               @      �?              G@      *@      @      @      @      @      @      @       @               @      @              �?       @       @              �?      �?             �D@      "@      D@      @      ;@      @      7@      @      6@      @      @      @      @      �?      �?      @               @      �?       @      2@              �?              @      �?      @                      �?      *@      �?      @              "@      �?      @               @      �?              �?       @              �?       @               @      �?             �B@      �?      3@              2@      �?       @              0@      �?       @      �?      ,@             @m@      k@     �a@     �d@     �[@     �Y@      <@      M@      �?     �J@               @      �?     �F@      �?      6@              "@      �?      *@      �?      @      �?                      @              "@              7@      ;@      @      @      @       @      @       @      �?       @                      �?               @       @              7@       @      7@                       @     �T@      F@     �T@     �E@     �N@      D@      (@      $@      �?      @              @      �?              &@      @      $@       @      @       @      @              �?       @               @      �?              @              �?      @              @      �?             �H@      >@      H@      :@      ;@      4@      ;@      0@      7@      0@      @       @      @      �?      �?      �?      �?                      �?      @                      �?      3@      ,@      2@      &@      (@      &@              "@      (@       @      @       @      @              @       @      @              �?       @      @              @              �?      @      �?      �?               @      @                      @      5@      @      5@      @              @      5@       @      4@       @      $@       @       @               @       @               @       @              $@              �?                      �?      �?      @      �?                      @      5@      @              @      5@                      �?      @@      P@      8@      P@      "@       @      �?      @              @      �?      �?      �?                      �?       @       @       @                       @      .@      L@      &@     �J@      "@     �J@      @      ,@      @      ,@              $@      @      @      �?      @              @      �?      �?              �?      �?               @              @              @     �C@       @     �A@       @      =@              0@       @      *@              @       @      @      �?      @              @      �?      @               @      �?      �?      �?                      �?      �?                      @      �?      @              @      �?               @              @      @      �?              @      @      @       @      @                       @              �?       @              W@     �I@      2@      7@      @      1@      @      1@              @      @      &@      �?              @      &@               @      @      "@      @      @      @                      @               @       @              (@      @      @      @      @      �?              �?      @              �?      @      �?      �?      �?                      �?              @      @             �R@      <@     �A@      9@      *@      1@      @      *@       @      *@       @       @       @      �?              �?       @                      �?              &@      �?              $@      @      @      @      @                      @      @              6@       @              @      6@      @      @      @      �?      @      �?                      @      @              2@             �C@      @       @      @      @              @      @      @              �?      @               @      �?      �?      �?                      �?      ?@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ	�tlhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B@D         J                    �?�4�O��?�           8�@               5                    �?r�=���?~            �h@                                  �?T �����?[             c@      =@                           �?�i�y�?$            �O@     *@                           �?`Ӹ����?            �F@      @������������������������       �                     6@      3@                            @���}<S�?             7@      @������������������������       �                     @      @	       
                 ���@�����H�?             2@       @������������������������       �                      @       @������������������������       �        
             0@      �?������������������������       �        
             2@                                    �?��Hg���?7            �V@      �?                           �?և���X�?             5@     0@                           �?���Q��?             4@                               `f�A@�q�q�?             (@     �?������������������������       �                     @      �?������������������������       �                     @                                  �5@      �?              @      �?������������������������       �                      @                                  �H@r�q��?             @     �?������������������������       �                     @     3@������������������������       �                     �?      C@������������������������       �                     �?      @                        ���@�~t��?*            @Q@        ������������������������       �        
             2@      �?       4                    �?��x_F-�?             �I@     ,@       3                 �|�=@j�q����?             I@              *                    �?      �?             B@     �?       %                   �:@���y4F�?             3@       @                         �&�)@�q�q�?             @        ������������������������       �                     �?        !       "                   �8@z�G�z�?             @      @������������������������       �                     @       @#       $                 �0@      �?              @       @������������������������       �                     �?      $@������������������������       �                     �?      @&       )                   @@8�Z$���?             *@       @'       (                 �|=@�q�q�?             @      @������������������������       �                      @      :@������������������������       �      �?             @       @������������������������       �                     @      �?+       .                 �|Y=@�t����?
             1@      &@,       -                  ��@      �?             @       @������������������������       �                      @       @������������������������       �                      @      �?/       2                    �?�θ�?             *@     @0       1                  s�@�z�G��?             $@       @������������������������       �                     @       @������������������������       �      �?             @      �?������������������������       �                     @      @������������������������       �                     ,@      P@������������������������       �                     �?      @6       C                    �?8�A�0��?#             F@      @7       <                 �|Y=@�LQ�1	�?             7@    �J@8       ;                 03�-@r�q��?
             (@      $@9       :                    &@�q�q�?             @      �?������������������������       �                     �?        ������������������������       �                      @      0@������������������������       �                     "@      @=       B                    �?�eP*L��?	             &@     �?>       ?                   @E@r�q��?             @      @������������������������       �                     @        @       A                 <3gH@�q�q�?             @       @������������������������       �                     �?        ������������������������       �                      @      1@������������������������       �                     @      &@D       I                     @؇���X�?             5@       E       H                 �̾w@�θ�?             *@     @F       G                    )@�C��2(�?
             &@        ������������������������       �                     �?      �?������������������������       �        	             $@      9@������������������������       �                      @       @������������������������       �                      @      �?K       �                    �?D����?C           �@      @L       m                    �?�BA����?f            `d@       @M       l                   �J@�7�QJW�?/            �R@     @N       [                     @v���a�?.            @R@       O       P                   �6@$�q-�?             J@      @������������������������       �        	             2@      �?Q       Z                   �*@�t����?             A@        R       S                   �'@�	j*D�?
             *@        ������������������������       �                      @        T       U                    :@���|���?             &@        ������������������������       �                      @        V       W                   �B@�<ݚ�?             "@       ������������������������       �                     @        X       Y                    D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     5@        \       k                    @�q�q�?             5@       ]       j                 @�"@�z�G��?             4@       ^       i                 `��!@և���X�?
             ,@       _       b                 ���@�q�q�?	             (@        `       a                 �|Y:@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        c       d                    4@և���X�?             @        ������������������������       �                      @        e       f                 @3�@z�G�z�?             @       ������������������������       �                     @        g       h                 �|Y>@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        n       �                 �D�H@��7��?7             V@       o       �                    @�{r٣��?'            �P@       p       q                    @JJ����?            �G@        ������������������������       �                     @        r       �                    �?�D����?             E@       s       �                    @\�Uo��?             C@       t       u                   �6@և���X�?            �A@        ������������������������       �                     @        v       }                     @     ��?             @@        w       x                   �7@      �?             (@        ������������������������       �                      @        y       |                    �?ףp=
�?             $@       z       {                    D@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ~                        �|Y=@�z�G��?             4@        ������������������������       �                     @        �       �                    �?���Q��?             .@        �       �                 ��1@�q�q�?             @01310,7������������������������       �                     @ 5,,Q
36������������������������       �                      @,7.25,,�       �                 `fV6@�<ݚ�?             "@ n)",fem������������������������       �                     �? oura Bo�       �                 ��T?@      �?              @Annie",������������������������       �                     @Pauline������������������������       �                     �? George ������������������������       �                     @nd, Mr. �       �                    �?      �?             @ an, Mr.������������������������       �                      @ghini, M������������������������       �                      @son, Mis�       �                 pfv2@p�ݯ��?
             3@ yer, Mr������������������������       �                     @8,,C
37�       �                    �?$�q-�?             *@ 077,7.2������������������������       �                      @ 03,211.�       �                 ��T?@z�G�z�?             @0125,,C������������������������       �                     @ ,7.775,������������������������       �                     �?7,227.52�       �                    #@�C��2(�?             6@ ,2653,1������������������������       �                     �? 2. 310�       �                 ���P@���N8�?             5@ ary Ali������������������������       �                     $@ky, Mr.�       �                 X�,@@�C��2(�?             &@ harles �       �                    �?�q�q�?             @  Master������������������������       �                     �?ss, Miss�       �                 ���d@      �?              @ atthew"������������������������       �                     �? a",fema������������������������       �                     �? st",mal������������������������       �                      @ Olof",m�       �                     �?PN��T'�?�            �u@ n Birge�       �                   �>@�j�'�=�?*            �P@ rjorie"�       �                   �<@r�q��?             8@ s. Hjal������������������������       �                     @.7,G6,S�       �                   �Q@��Q��?             4@,S
397,�       �                   @E@�E��ӭ�?             2@398,0,2�       �                 03:@d}h���?
             ,@ 2,"Pain������������������������       �                      @ Mrs. Wi�       �                 03k:@      �?             @ ,"Niska������������������������       �                     �?2,0,3,"A�       �                 �|�?@���Q��?             @la, Mis�       �                 `fF<@      �?             @ ainen, ������������������������       �                      @405,0,3�       �                 �|Y=@      �?              @ 
406,0,������������������������       �                     �? idegren������������������������       �                     �? 1,2,"Ri������������������������       �                     �?09,0,3,�       �                    K@      �?             @775,,S
�       �                   @G@�q�q�?             @411,0,3������������������������       �      �?              @ "Hart, ������������������������       �                     �?iss. Da������������������������       �                     �?Mr. Alf������������������������       �                      @ Johan J�       �                 �|�<@��s����?             E@ ek, Mrs������������������������       �                     @ S
417,1�       �                    �?�ݜ�?            �C@le,34,1�       �                   �E@4?,R��?             B@female,�       �                  x#J@�E��ӭ�?             2@male,30������������������������       �                     "@ale,10,0�       �                 �|Y>@X�<ݚ�?             "@ ,0,0,34������������������������       �                      @ A/5. 13�       �                 `f�K@����X�?             @ 5082,7.�       �                 `�iJ@�q�q�?             @ aria Br������������������������       �                     �?. Vikto������������������������       �                      @, Mr. P������������������������       �                     @Mrs. Cha������������������������       �        	             2@,1,2,"P������������������������       �                     @ Marshal�       �                    '@�W�{�5�?�            �q@ s",male�       �                     @��H�}�?             9@ mbisky)������������������������       �                     @strom-S�       �                 ���A@      �?
             2@52,S
43�       �                    @ףp=
�?             $@ ,female������������������������       �                     �?der (Ali������������������������       �                     "@3,"Kalli������������������������       �                      @ 5,,S
43�       �                 �?�@0Oex�I�?�            @p@ E44,S
4�       �                     @p� V�?=            �Y@ 20,B96 ������������������������       �                     @emale,21�       �                    ?@@��8��?9             X@(Emily �       �                   �8@@�z�G�?.             T@ Mr. Mar�       �                    7@ ���J��?            �C@ Mr. Jo������������������������       �                     ?@1,1,2,"�       �                 `fF@      �?              @ 1,F.C.C�       �                 �&b@�q�q�?             @ 5769,9.������������������������       �                      @76,7.77������������������������       �                     �?30434,13������������������������       �                     @,65306,������������������������       �                    �D@,33638,8�       �                 �&B@      �?             0@female,������������������������       �        
             .@r",male������������������������       �                     �?herine"�                          �?P��-�?h            �c@thur Go�       �                     @0�I��8�?T             _@ Edwy Ar�       �                    F@dP-���?!            �G@r. Ingv�       �                   @D@������?            �B@an, Mr.�       �                   �3@�#-���?            �A@1,1,"Go�       �                   �(@ȵHPS!�?             :@ 55,0,3,�       �                   �5@$�q-�?             *@ "Jalsev�       �                    &@r�q��?             @ t, Mr. ������������������������       �                     �?nyon, Mr������������������������       �                     @ 459,1,2������������������������       �                     @S
460,0,�       �                 �|�<@8�Z$���?
             *@ 1,"Ande������������������������       �                     @orley, �       �                   �A@�q�q�?             @ Arthur�       �                 �|�=@�q�q�?             @ acob Ch������������������������       �                     �?Simon",m�       �                    @@      �?              @ Estansl������������������������       �                     �?bell, Mr������������������������       �                     �? Montgo������������������������       �                     @ ames",m������������������������       �                     "@ rbara",������������������������       �      �?              @ r",male������������������������       �                     $@0,31508�                         @@@؇���X�?3            @S@th)",fe�       
                �|Y>@���*�?&             N@n S (Ma�                       �!&B@�t����?!            �I@917,D,C�       �                   �1@�8��8��?             H@ ,9.8375������������������������       �                     $@5,52,A1�       �                   �2@�KM�]�?             C@ 1,,S
47������������������������       �                     �?8,,S
479�       �                 ��) @�L���?            �B@ 8,,S
48������������������������       �                     4@.2875,,S�                       @3�!@@�0�!��?             1@ 144,46.�       �                 pf� @�q�q�?             @ ,0,2398������������������������       �                     �?5 3594,                       �|Y<@      �?              @ 34,9.58������������������������       �                     �?        ������������������������       �                     �?                                �<@@4և���?             ,@       ������������������������       �                     &@                              �|Y=@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @              	                   ;@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                �?@X�<ݚ�?             "@        ������������������������       �                     @                              ��I @�q�q�?             @       ������������������������       ����Q��?             @        ������������������������       �                     �?        ������������������������       �                     1@        ������������������������       �                    �@@        �t�bh�h*h-K ��h/��R�(KMKK��h]�B       �{@     �p@      X@     @Y@     �Q@     �T@       @     �N@       @     �E@              6@       @      5@              @       @      0@       @                      0@              2@      Q@      6@      "@      (@       @      (@      @      @              @      @              @      @       @              �?      @              @      �?              �?             �M@      $@      2@             �D@      $@     �D@      "@      ;@      "@      .@      @      @       @              �?      @      �?      @              �?      �?      �?                      �?      &@       @      @       @       @               @       @      @              (@      @       @       @       @                       @      $@      @      @      @      @              @      @      @              ,@                      �?      :@      2@       @      .@       @      $@       @      �?              �?       @                      "@      @      @      �?      @              @      �?       @      �?                       @      @              2@      @      $@      @      $@      �?              �?      $@                       @       @             �u@     `d@      J@     �[@      *@      O@      &@      O@      @      H@              2@      @      >@      @      "@               @      @      @       @               @      @              @       @      �?       @                      �?              5@      @      ,@      @      ,@      @       @      @       @      �?      @              @      �?              @      @       @              �?      @              @      �?      �?      �?                      �?       @                      @      �?               @             �C@     �H@     �B@      =@      9@      6@              @      9@      1@      7@      .@      4@      .@      @              1@      .@      @      "@       @              �?      "@      �?      @              @      �?                      @      ,@      @      @              "@      @       @      @              @       @              @       @              �?      @      �?      @                      �?      @               @       @               @       @              (@      @              @      (@      �?       @              @      �?      @                      �?       @      4@      �?              �?      4@              $@      �?      $@      �?       @              �?      �?      �?      �?                      �?               @     �r@      J@     �G@      3@      *@      &@              @      *@      @      *@      @      &@      @       @              @      @              �?      @       @      @      �?       @              �?      �?      �?                      �?              �?       @       @      �?       @      �?      �?              �?      �?                       @      A@       @              @      A@      @      ?@      @      *@      @      "@              @      @       @               @      @       @      �?              �?       @                      @      2@              @             �o@     �@@      "@      0@              @      "@      "@      �?      "@      �?                      "@       @             `n@      1@     @Y@       @      @             �W@       @     �S@      �?      C@      �?      ?@              @      �?       @      �?       @                      �?      @             �D@              .@      �?      .@                      �?     �a@      .@     @[@      .@     �E@      @     �@@      @      @@      @      7@      @      (@      �?      @      �?              �?      @              @              &@       @      @              @       @      �?       @              �?      �?      �?      �?                      �?      @              "@              �?      �?      $@             �P@      &@     �H@      &@     �F@      @      F@      @      $@              A@      @              �?      A@      @      4@              ,@      @      �?       @              �?      �?      �?              �?      �?              *@      �?      &@               @      �?              �?       @              �?       @               @      �?              @      @              @      @       @      @       @      �?              1@             �@@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�ޡhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM%huh*h-K ��h/��R�(KM%��h|�B@I         �                 `f~I@�t����?�           8�@ X         S                    �?�����2�?�           h�@                                ��@V���#�?~            �g@ pñX                          �|Y:@�IєX�?             1@5.3"}�?������������������������       �                     &@ will be                        �&�@r�q��?             @ turns
 ������������������������       �                     �?essions ������������������������       �                     @ach valu	                            @�.�8�?q            �e@      �?
                        ���*@�L#���?/            �P@      @                        `f�)@      �?             8@       @                          �J@$�q-�?             *@      @������������������������       �                     (@        ������������������������       �                     �?       @                          �B@"pc�
�?	             &@                                  :@�����H�?             "@      @                           �?�q�q�?             @      �?������������������������       �                     �?        ������������������������       �                      @      �?������������������������       �                     @                                   D@      �?              @      �?������������������������       �                     �?     3@������������������������       �                     �?      C@                           E@ qP��B�?            �E@     @������������������������       �                     ?@                                    �?�8��8��?             (@      �?������������������������       �                     @     ,@                           �?r�q��?             @        ������������������������       �                     �?     �?������������������������       �                     @       @       &                    @�k��V��?B            �Z@                %                    �?؇���X�?             ,@       !       $                    @      �?              @      0@"       #                 ��0@      �?             @      "@������������������������       �                      @     @������������������������       �                      @     �?������������������������       �                     @     @������������������������       �                     @     0@'       D                 03�1@�+Fi��?;             W@     *@(       =                 �?�-@�ݜ����?'            �M@     @)       ,                 �̌@�&!��?            �E@       @*       +                   �2@�z�G��?             $@        ������������������������       �                     @      @������������������������       �                     @      �?-       .                   �1@:ɨ��?            �@@      @������������������������       �                     @      �?/       <                    �?PN��T'�?             ;@     @0       1                 `�X!@���y4F�?             3@      �?������������������������       �                     @       @2       7                   �9@����X�?	             ,@     �?3       6                    4@      �?              @      �?4       5                    �?�q�q�?             @      �?������������������������       �                      @     �?������������������������       �                     �?     �?������������������������       �                     @      4@8       9                    �?      �?             @      (@������������������������       �                     �?      @:       ;                    A@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @      @������������������������       �                      @      �?>       ?                   �0@      �?
             0@      @������������������������       �                     �?        @       C                   �;@��S�ۿ?	             .@        A       B                    �?�q�q�?             @       @������������������������       �                     �?      �?������������������������       �                      @      �?������������������������       �                     (@        E       H                    @"pc�
�?            �@@       F       G                    �?�����?             5@        ������������������������       �                      @        ������������������������       �                     3@        I       J                 0C�7@�q�q�?             (@        ������������������������       �                     �?        K       L                    �?���!pc�?             &@        ������������������������       �                     @        M       N                    @      �?              @        ������������������������       �                      @        O       R                    @      �?             @       P       Q                   @C@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        T       m                 �?�@б΅t�?           �x@        U       l                    �?�wY;��?X             a@       V       k                 �Yu@     x�?S             `@       W       b                    �?���F6��?B            �X@        X       Y                 ���@�ݜ�?            �C@        ������������������������       �        	             .@        Z       [                   �6@�q�q�?             8@        ������������������������       �                      @        \       ]                  ��@��2(&�?             6@        ������������������������       �                     "@        ^       _                 �|Y=@�θ�?	             *@        ������������������������       �                     �?        `       a                 X��A@r�q��?             (@       ������������������������       �z�G�z�?             $@        ������������������������       �                      @        c       d                    7@(;L]n�?)             N@        ������������������������       �                     3@        e       j                 ��L@������?            �D@       f       g                 ���@�(\����?             D@        ������������������������       �                     5@        h       i                 ���@�}�+r��?             3@        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     �?        ������������������������       �                     =@        ������������������������       �                      @        n       �                     �?|;�c� �?�            pp@        o       t                 �|�<@�q�q�?              H@        p       q                   �;@؇���X�?             @        ������������������������       �                      @        r       s                 `f�D@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        u       �                    �?���?            �D@       v       �                  �>@�d�����?             C@       w       �                    K@���Q��?             9@       x       �                   �G@���Q��?
             .@       y       ~                    �?���Q��?             $@        z       {                 `f&;@      �?             @        ������������������������       �                      @        |       }                 �|�=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @               �                 03k:@      �?             @        �       �                   �D@      �?              @        ������������������������       �                     �?1.275,,S������������������������       �                     �?v�X  ������������������������       �                      @%��X  ������������������������       �                     @8?�X  �       �                 ���=@ףp=
�?             $@emale,4������������������������       �                     "@female,1������������������������       �                     �?(Mary Hi������������������������       �        	             *@ Mr. Pet������������������������       �                     @�l�X  �       �                    �?��ݼ��?�            �j@:�X  �       �                     @�r����?W            �`@ en, Mr.�       �                    �? "��u�?              I@ C�X  ������������������������       �                     �?ft, Mrs.�       �                    �?��<D�m�?            �H@7466,25�       �                   �*@      �?             H@,female�       �                 `fF)@l��\��?             A@ male,24������������������������       �                     $@��X  �       �                 �|�<@      �?             8@ male,27������������������������       �                     *@hington �       �                   �F@���!pc�?             &@van Mel�       �                 �|�=@      �?             @ �X  ������������������������       �                     �?���X  �       �                    B@���Q��?             @ ckwith,������������������������       �                      @cU�X  ������������������������       ��q�q�?             @0,695,5,������������������������       �                     @#E�X  ������������������������       �                     ,@y)",fema������������������������       �                     �?"��X  �       �                    �?@�0�!��?7            @U@ r. Alfr������������������������       �                     @Mr. Nede�       �                 @3�@����!�?4            �T@ ��X  �       �                    :@�eP*L��?             &@  (Lily ������������������������       �                     @1,2,"She�       �                   �?@����X�?             @ ��X  ������������������������       �                      @8958,,S
�       �                   �A@���Q��?             @ ,10.516������������������������       ��q�q�?             @,C.A./SO������������������������       �      �?              @�?�X  �       �                    )@D��\��?-            �Q@ ret Nor������������������������       �                     �?Rev. Juo�       �                 �|Y=@������?,            �Q@ aret Ed�       �                 ��Y @��a�n`�?             ?@ ��X  �       �                   �3@      �?              @ 90,1,1,������������������������       �                     @��X  ������������������������       �                     @^� �0�u �       �                 `�X#@�㙢�c�?             7@^�X  �       �                 ���"@���y4F�?             3@��X  �       �                 @�!@�r����?
             .@       �       �                 pf� @�<ݚ�?             "@        ������������������������       �                      @�$�X  �       �                    8@����X�?             @��X  ������������������������       �                     @i��X  ������������������������       �                      @        ������������������������       �                     @I|�X  �       �                   �<@      �?             @       ������������������������       �                      @��X  ������������������������       �                      @        ������������������������       �                     @�%�X  �       �                   �?@�7��?            �C@M�X  �       �                 ��) @���}<S�?             7@       ������������������������       �                     ,@0^�X  �       �                 �|�=@�<ݚ�?             "@q�X  �       �                 pf� @      �?              @ &�X  ������������������������       �                     �?���X  ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             0@��X  �       �                    �?�z�G��?5             T@ �X  �       �                 �2@�n_Y�K�?             *@       �       �                 �|�;@�����H�?             "@       �       �                 �&�)@      �?             @ �X  ������������������������       �                      @N��X  �       �                    �?      �?              @ p�X  ������������������������       �                     �?        ������������������������       �                     �?>9�X  ������������������������       �                     @        ������������������������       �                     @���X  �       �                    �?���}D�?-            �P@ @�X  �       �                    �? ��WV�?             :@ ��X  ������������������������       �                     @        �       �                    6@�nkK�?             7@        ������������������������       �                     �?        ������������������������       �                     6@        �       �                    @��]�T��?            �D@3�X  �       �                    �?\�Uo��?             C@ ��X  ������������������������       �                      @G��X  �       �                    @�q�q�?             B@4�X  �       �                 03{3@�q�����?             9@        �       �                     @z�G�z�?             $@ l�X  �       �                    *@z�G�z�?             @ ��X  ������������������������       �                     �?��X  ������������������������       �                     @S3�X  �       �                   �5@z�G�z�?             @C�X  ������������������������       �                     @w��X  ������������������������       �                     �?        �       �                 �̌4@�q�q�?             .@ .�X  ������������������������       �                     @        �       �                    �?�q�q�?             (@��X  �       �                    :@�z�G��?             $@       �       �                     @      �?             @        ������������������������       �                      @        �       �                    +@      �?              @ ��X  ������������������������       �                     �?        ������������������������       �                     �?�.�X  ������������������������       �                     @        ������������������������       �                      @        �       �                    �?"pc�
�?             &@        ������������������������       �                     @���X  �       �                 pf�C@�q�q�?             @        �       �                    @�q�q�?             @        ������������������������       �                      @8s�X  ������������������������       �                     �?h��X  ������������������������       �                     @        ������������������������       �                     @        �       �                    �?ƆQ����?P            �^@��X  �       �                  "�b@pY���D�?0            �S@       ������������������������       �        %            �M@        �       �                    �?ףp=
�?             4@L�X  ������������������������       �                     $@        �       �                    $@z�G�z�?             $@ \�X  ������������������������       �                      @�)�X  ������������������������       �                      @        �                           @�&!��?             �E@       �                          �?p�ݯ��?             C@��X  �                           �?b�2�tk�?             B@       �       	                �UwR@���Q��?            �A@ �X  �                          �?�<ݚ�?             2@                                  �?���Q��?             @        ������������������������       �                      @                              ��UO@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                �C@$�q-�?             *@        ������������������������       �                     @                                 F@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        
                         �?j���� �?             1@                                 �?      �?              @                                �?؇���X�?             @                                �9@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?                                 �?X�<ݚ�?             "@                                �?z�G�z�?             @                              �̾w@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                 �?      �?             @                                =@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @              $                p�O@���Q��?             @              #                   >@      �?             @       !      "                   ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �t�b�[     h�h*h-K ��h/��R�(KM%KK��h]�BP       �z@     �q@     �x@      h@      O@      `@      �?      0@              &@      �?      @      �?                      @     �N@      \@      @     �O@      @      5@      �?      (@              (@      �?               @      "@      �?       @      �?       @      �?                       @              @      �?      �?      �?                      �?      �?      E@              ?@      �?      &@              @      �?      @      �?                      @     �L@     �H@       @      (@       @      @       @       @               @       @                      @              @     �K@     �B@      <@      ?@      :@      1@      @      @      @                      @      7@      $@              @      7@      @      .@      @      @              $@      @      @      �?       @      �?       @                      �?      @              @      @      �?               @      @              @       @               @               @      ,@      �?              �?      ,@      �?       @      �?                       @              (@      ;@      @      3@       @               @      3@               @      @              �?       @      @      @              @      @       @              @      @       @      @              @       @              �?             �t@     @P@      `@      @     @^@      @      W@      @      A@      @      .@              3@      @               @      3@      @      "@              $@      @              �?      $@       @       @       @       @              M@       @      3@             �C@       @     �C@      �?      5@              2@      �?              �?      2@                      �?      =@               @             �i@      M@      @@      0@      �?      @               @      �?      @              @      �?              ?@      $@      <@      $@      .@      $@      @      "@      @      @      @      @               @      @      �?              �?      @              @      �?      �?      �?              �?      �?               @                      @      "@      �?      "@                      �?      *@              @             �e@      E@     @]@      2@     �G@      @      �?              G@      @     �F@      @      ?@      @      $@              5@      @      *@               @      @      @      @              �?      @       @       @              �?       @      @              ,@              �?             �Q@      .@      @             �P@      .@      @      @      @               @      @               @       @      @      �?       @      �?      �?     �N@      $@              �?     �N@      "@      8@      @      @      @              @      @              3@      @      .@      @      *@       @      @       @       @              @       @      @                       @      @               @       @       @                       @      @             �B@       @      5@       @      ,@              @       @      @      �?              �?      @                      �?      0@              L@      8@      @       @      �?       @      �?      @               @      �?      �?      �?                      �?              @      @             �I@      0@      9@      �?      @              6@      �?              �?      6@              :@      .@      7@      .@       @              5@      .@      (@      *@       @       @      �?      @      �?                      @      �?      @              @      �?              $@      @      @              @      @      @      @      �?      @               @      �?      �?              �?      �?              @                       @      "@       @      @              @       @      �?       @               @      �?              @              @              <@     �W@       @     @S@             �M@       @      2@              $@       @       @       @                       @      :@      1@      8@      ,@      6@      ,@      5@      ,@      ,@      @       @      @               @       @      �?       @                      �?      (@      �?      @              @      �?              �?      @              @      $@       @      @      �?      @      �?       @      �?                       @              @      �?              @      @      @      �?      �?      �?      �?                      �?      @              �?      @      �?      �?              �?      �?                       @      �?               @               @      @      �?      @      �?      �?              �?      �?                       @      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJQY%hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtK�huh*h-K ��h/��R�(KK���h|�B�?                             @��ϙLq�?�           8�@      0@       	                    @     ��?             @@     @                           @��.k���?             1@     =@                           �?ףp=
�?             $@      *@                             @      �?              @      �?������������������������       �                     �?      0@������������������������       �                     �?      "@������������������������       �                      @        ������������������������       �                     @0(Y�X  
                           �?��S�ۿ?
             .@"Y�X  ������������������������       �                     $@�2Y�X                             @z�G�z�?             @ +Y�X  ������������������������       �                     @�2Y�X                             �?      �?              @ 0Y�X  ������������������������       �                     �?        ������������������������       �                     �?0$Y�X         �                 `fK@�ĸۦ��?�           8�@     �?       Q                    �?��J��?r           @�@               "                     @Z�2�t��?h            �d@      �?       !                    �?0)RH'�?(            @Q@                                 �*@�q�q��?             H@      �?                           B@���Q��?             4@     3@                          �9@      �?	             0@      C@                          �'@z�G�z�?             @      @������������������������       �                     �?        ������������������������       �                     @      �?������������������������       �                     &@     ,@������������������������       �                     @                                ���;@ �Cc}�?             <@     �?������������������������       �                     6@       @                         X��C@      �?             @       ������������������������       �                     @       ������������������������       �                     @      @������������������������       �                     5@        #       0                 pF @�W*��?@            @X@      �?$       /                    �?��hJ,�?             A@     @%       .                 X��B@<���D�?            �@@      @&       '                   �6@     ��?             @@        ������������������������       �                     .@        (       )                   �8@@�0�!��?             1@        ������������������������       �                      @      @*       -                 ���@��S�ۿ?             .@        +       ,                 �Y�@      �?             @      @������������������������       �                     @       @������������������������       �                     �?      �?������������������������       �        	             &@        ������������������������       �                     �?      @������������������������       �                     �?      @1       N                 03�7@����X�?+            �O@       2       K                    �?�D����?             E@     �?3       F                    �?p�ݯ��?             C@     @4       ?                 ��.@     ��?             @@     &@5       >                    �?�J�4�?             9@       6       ;                 �&�%@������?             1@     (@7       :                 `��!@ףp=
�?             $@      @8       9                 `�X!@      �?             @      @������������������������       �                     @      �?������������������������       �                     �?        ������������������������       �                     @      �?<       =                 ���*@և���X�?             @      $@������������������������       �                     @       @������������������������       �                     @       @������������������������       �                      @      @@       A                    �?؇���X�?             @       @������������������������       �                     @      �?B       C                 03�1@      �?             @      �?������������������������       �                      @      @D       E                    �?      �?              @      @������������������������       �                     �?      �?������������������������       �                     �?      @G       J                    @�q�q�?             @      @H       I                   �4@���Q��?             @      @������������������������       �                      @       @������������������������       �                     @        ������������������������       �                     �?        L       M                 �|Y=@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        O       P                    �?���N8�?             5@        ������������������������       �                     �?        ������������������������       �                     4@        R       �                   �J@T�1!�}�?
            z@       S       \                   �2@      �?�            �x@        T       [                 �&@������?             B@        U       V                    �?�X�<ݺ?             2@       ������������������������       �                     $@        W       Z                    �?      �?              @        X       Y                  �K"@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     2@        ]       x                     �?4�<����?�            @v@        ^       e                 �|�<@��J�fj�?            �B@        _       `                    7@      �?              @        ������������������������       �                     �?        a       b                 `f�D@؇���X�?             @       ������������������������       �                     @        c       d                 ��I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        f       w                   �G@J�8���?             =@       g       r                 �TA@@l��
I��?             ;@       h       m                 ���=@j���� �?             1@       i       l                 ��";@"pc�
�?
             &@       j       k                 ��:@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        n       o                  �>@r�q��?             @        ������������������������       �                     @        p       q                  �>@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        s       t                   �C@ףp=
�?             $@       ������������������������       �                     @        u       v                    �?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        y       �                    �?0�\>��?�            �s@       z       �                   @E@�u����?�             q@       {       �                    �?Ǖi�7�?�            0p@       |       �                     @X�EQ]N�?�             p@        }       ~                    �?���c���?             J@        ������������������������       �                     @               �                   @D@؇���X�?            �H@       �       �                 `fF)@�����H�?            �F@        �       �                    5@���7�?             6@        ������������������������       �                     �?        ������������������������       �                     5@        �       �                 �|�<@�㙢�c�?             7@        ������������������������       �                      @        �       �                   �3@������?             .@       �       �                   �A@�	j*D�?             *@       �       �                    @@      �?              @       �       �                 �|�=@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �      �?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �      �?             @        �       �                 �Y�@�"�_*d�?�            �i@        �       �                   �8@���y4F�?             C@        �       �                   �3@���|���?             &@        ������������������������       �                     @        �       �                    5@      �?              @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ���@ 7���B�?             ;@       ������������������������       �                     6@       ������������������������       �z�G�z�?             @        �       �                 �?�@4և����?k             e@       �       �                 �?$@x��B�R�?9            �V@        �       �                    ;@�8��8��?             B@        ������������������������       �                     *@        �       �                  s�@�LQ�1	�?             7@        ������������������������       �                     @        �       �                    �?     ��?             0@       �       �                 �|Y=@"pc�
�?	             &@        ������������������������       �                     �?        �       �                 X��A@ףp=
�?             $@       ������������������������       ������H�?             "@       ������������������������       �                     �?        �       �                 �|Y>@z�G�z�?             @        ������������������������       �      �?              @        ������������������������       �                     @        ������������������������       �                    �K@        �       �                    �?� ���?2            @S@        ������������������������       �                     @        �       �                   @C@�MI8d�?/            �R@       �       �                   �3@؇���X�?,            �Q@        ������������������������       ����Q��?             @        �       �                 ��) @�?�<��?*            @P@       �       �                   �>@��(\���?             D@       ������������������������       �                     =@        �       �                   �@@���!pc�?             &@       �       �                   �?@      �?             @        ������������������������       �                     �?        ������������������������       ����Q��?             @        ������������������������       �                     @        �       �                 �|�>@z�G�z�?             9@       �       �                   �8@      �?             4@        ������������������������       �                     @        �       �                 0S%"@     ��?             0@        �       �                 �|Y<@���Q��?             @        ������������������������       �                      @        �       �                 pf� @�q�q�?             @        ������������������������       �                     �?       ������������������������       �                      @       �       �                   �<@"pc�
�?             &@        ������������������������       �                     @        �       �                 �|Y=@���Q��?             @        �       �                 ���"@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   @D@      �?             @       �       �                 ��	0@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?       ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     .@        �       �                 ��.@`Ӹ����?            �F@        �       �                    �?r�q��?	             (@       �       �                     @�C��2(�?             &@        ������������������������       �                     �?       �       �                    5@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@       ������������������������       �                     �?        ������������������������       �                    �@@        ������������������������       �                     :@        �       �                    �?�"�q��?A            �W@       �       �                    �?�}�+r��?'            �L@       ������������������������       �                     =@       �       �                    @ �Cc}�?             <@       ������������������������       �                     9@        ������������������������       �                     @       �       �                    �?p�ݯ��?             C@       �       �                 X�,@@��Q��?             4@       �       �                  �}S@      �?             $@        ������������������������       �                     @        �       �                    �?r�q��?             @       ������������������������       �                     @        �       �                   �5@      �?              @        ������������������������       �                     �?       ������������������������       �                     �?       �       �                    �?z�G�z�?             $@       �       �                   @H@�����H�?             "@       ������������������������       �                     @        �       �                   �T@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                     @b�2�tk�?             2@       �       �                     �?      �?	             (@       �       �                 �|Y>@�eP*L��?             &@        ������������������������       �                     �?       �       �                    �?���Q��?             $@       �       �                 03�U@      �?              @       �       �                    C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?       �       �                    @r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KK�KK��h]�B�       �|@     �o@      "@      7@       @      "@      �?      "@      �?      �?      �?                      �?               @      @              �?      ,@              $@      �?      @              @      �?      �?      �?                      �?     �{@      m@     �z@     @c@     �N@     @Z@      &@      M@      &@     �B@       @      (@      @      (@      @      �?              �?      @                      &@      @              @      9@              6@      @      @              @      @                      5@      I@     �G@      @      =@      @      =@      @      =@              .@      @      ,@       @              �?      ,@      �?      @              @      �?                      &@      �?              �?             �F@      2@      9@      1@      8@      ,@      6@      $@      5@      @      *@      @      "@      �?      @      �?      @                      �?      @              @      @              @      @               @              �?      @              @      �?      @               @      �?      �?      �?                      �?       @      @       @      @       @                      @              �?      �?      @              @      �?              4@      �?              �?      4@             w@     �H@     pu@     �H@     �A@      �?      1@      �?      $@              @      �?      @      �?      @                      �?      @              2@             @s@      H@      5@      0@       @      @      �?              �?      @              @      �?      �?      �?                      �?      3@      $@      3@       @      $@      @      "@       @      @       @      @                       @      @              �?      @              @      �?       @      �?                       @      "@      �?      @              @      �?      @                      �?               @     �q@      @@     �n@      >@     �l@      >@     �l@      >@     �F@      @      @              E@      @      D@      @      5@      �?              �?      5@              3@      @       @              &@      @      "@      @      @      @      @      �?              �?      @              �?      @      @               @               @       @     �f@      7@      >@       @      @      @      @              �?      @      �?       @               @      �?                      @      :@      �?      6@              @      �?      c@      .@      V@      @     �@@      @      *@              4@      @      @              *@      @      "@       @              �?      "@      �?       @      �?      �?              @      �?      �?      �?      @             �K@             @P@      (@      @              O@      (@      N@      $@      @       @     �L@       @     �B@      @      =@               @      @      @      @              �?      @       @      @              4@      @      .@      @      @              &@      @       @      @               @       @      �?              �?       @              "@       @      @              @       @      �?       @      �?                       @       @              @               @       @      �?       @               @      �?              �?              �?              .@             �E@       @      $@       @      $@      �?      �?              "@      �?              �?      "@                      �?     �@@              :@              1@     �S@      @      K@              =@      @      9@              9@      @              ,@      8@      @      *@      @      @              @      @      �?      @              �?      �?      �?                      �?       @       @      �?       @              @      �?       @               @      �?              �?              @      &@      @      @      @      @      �?              @      @       @      @       @      �?              �?       @                      @       @              �?              �?      @              @      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ��fbhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM5huh*h-K ��h/��R�(KM5��h|�B@M         F                    �?�u����?�           8�@    tati                           �?sYi9��?O            `a@ ��X                              @\#r��?"            �N@    �Q@                          �H@��<b�ƥ?             G@     �?������������������������       �                     E@                                   J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        	                           �?�q�q�?
             .@     =@
                           �?X�Cc�?	             ,@      ,@                        �&�)@և���X�?             @      @������������������������       �                     @        ������������������������       �                     @      $@                        `�@1@����X�?             @     �?                           @      �?             @      @������������������������       �                      @      @������������������������       �                      @      �?������������������������       �                     @      @������������������������       �                     �?      @       E                 �U�X@�θ�?-            �S@     �?       D                  �	U@��R[s�?*            �Q@     �?       C                    �?��ga�=�?(            �P@     �?       <                 ��<J@�'�`d�?'            �P@              9                    �?&y�X���?#             M@              6                    �?r�����?             �J@              5                 p�i@@��k=.��?            �G@     @       2                   `A@�I�w�"�?             C@      @       1                 �|�=@"pc�
�?            �@@      @                             �?d}h���?             <@                                0C�<@      �?              @       @������������������������       �                     �?      >@������������������������       �                     �?      @!       (                    ;@���B���?             :@      @"       '                 ���@�8��8��?             (@       #       $                 ��y@؇���X�?             @      @������������������������       �                     �?      @%       &                   �7@r�q��?             @      @������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @      @)       *                 �|Y=@����X�?	             ,@      @������������������������       �                     �?      �?+       ,                     @�θ�?             *@      @������������������������       �                     �?       @-       0                   @@      �?             (@       .       /                 ���@      �?              @        ������������������������       �                     �?       @������������������������       �և���X�?             @      �?������������������������       �                     @      8@������������������������       �                     @       @3       4                      @���Q��?             @      @������������������������       �                     @        ������������������������       �                      @      .@������������������������       �                     "@      *@7       8                 �&�)@r�q��?             @      @������������������������       �                     �?      @������������������������       �                     @      @:       ;                ��k/@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        =       B                 ���Q@      �?              @    @S@>       A                    �?      �?             @      @?       @                    F@      �?              @      ,@������������������������       �                     �?      @������������������������       �                     �?      �?������������������������       �                      @      �?������������������������       �                     @      @������������������������       �                     �?      @������������������������       �                     @      �?������������������������       �                      @      @G                          �?��s�ɝ�?t           ��@      @H       �                    �?>4և���?"            |@     @I       z                    �?������?�            �w@       @J       g                   �9@z�G�z�?2            �R@        K       `                   �6@�û��|�?             7@       L       _                 8#B2@������?             1@       M       N                   �1@���|���?
             &@        ������������������������       �                     �?        O       X                   �4@���Q��?	             $@       P       Q                    �?      �?             @        ������������������������       �                     �?        R       W                    3@���Q��?             @       S       T                 P��@      �?             @        ������������������������       �                     �?        U       V                 ��!@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        Y       Z                     @      �?             @        ������������������������       �                     �?        [       \                    �?�q�q�?             @        ������������������������       �                     �?        ]       ^                 pF�!@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        a       b                     @r�q��?             @        ������������������������       �                     �?        c       f                    8@z�G�z�?             @       d       e                 @3�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @       ������������������������       �                      @       h       i                    �?ȵHPS!�?!             J@        ������������������������       �                     $@       j       w                     @؇���X�?             E@       k       n                 `f&'@ >�֕�?            �A@        l       m                   �E@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        o       p                     �?�g�y��?             ?@        ������������������������       �                     *@        q       r                   �B@�X�<ݺ?             2@       ������������������������       �                     "@        s       v                   �*@�����H�?             "@        t       u                    D@      �?             @        ������������������������       �                     �?       ������������������������       �                     @        ������������������������       �                     @        x       y                 �|�;@և���X�?             @        ������������������������       �                     @       ������������������������       �                     @       {       �                 ��$:@�Qb��?�            �r@       |       �                   @@@������?�            0p@       }       �                   �>@$�3c�s�?v            �g@       ~       �                 @3�@��I�� �?o            `f@              �                 �|Y=@��<D�m�?;            �X@        �       �                 ��@      �?             D@       �       �                  ��@z�G�z�?             9@01310,7�       �                    �?�C��2(�?             6@ 5,,Q
36������������������������       �                     �?,7.25,,�       �                    7@�����?             5@n)",fem������������������������       �                     (@ oura Bo�       �                 ���@�<ݚ�?             "@ Annie",�       �                 �&b@�q�q�?             @ Pauline������������������������       �                     �? George ������������������������       �                      @nd, Mr. ������������������������       �                     @ an, Mr.������������������������       �                     @ghini, M������������������������       �                     .@son, Mis�       �                 �|�=@ _�@�Y�?             M@yer, Mr�       �                     @@3����?             K@ 8,,C
37������������������������       �                     &@ 077,7.2�       �                 ��@ qP��B�?            �E@03,211.������������������������       �                     6@0125,,C�       �                 �Y5@���N8�?
             5@ ,7.775,������������������������       �z�G�z�?             @7,227.52������������������������       �                     0@ ,2653,1������������������������       �                     @ 2. 310�       �                   �3@�
��P�?4            @T@ ary Ali�       �                   �2@�d�����?             3@ky, Mr.�       �                 ��Y @ףp=
�?             $@ harles �       �                    1@      �?              @  Master������������������������       �                     �?ss, Miss������������������������       �                     �? atthew"������������������������       �                      @ a",fema�       �                 ���$@X�<ݚ�?             "@st",mal�       �                 0S5 @����X�?             @ Olof",m������������������������       ��q�q�?             @ n Birge������������������������       �                     @ rjorie"������������������������       �                      @ s. Hjal�       �                    �?��a�n`�?(             O@ .7,G6,S������������������������       �                     �?,S
397,�       �                 ��) @\#r��?'            �N@ 398,0,2������������������������       �                     6@ 2,"Pain�       �                    :@8�Z$���?            �C@ Mrs. Wi������������������������       �                     .@ ,"Niska�       �                     @      �?             8@ ,0,3,"A�       �                 �|Y<@�8��8��?             (@ la, Mis������������������������       �                     @ ainen, �       �                     �?؇���X�?             @ 405,0,3������������������������       �                      @ 
406,0,�       �                 �|�=@z�G�z�?             @ idegren������������������������       �                     �? 1,2,"Ri������������������������       �                     @09,0,3,�       �                 0S%"@�q�q�?             (@ 775,,S
�       �                 pf� @z�G�z�?             @ 411,0,3������������������������       �                      @ "Hart, �       �                 �|Y<@�q�q�?             @ iss. Da������������������������       �                      @Mr. Alf������������������������       �                     �? Johan J�       �                 �|�=@؇���X�?             @ek, Mrs������������������������       �                     @ S
417,1������������������������       �                     �?le,34,1�       �                 �&B@X�<ݚ�?             "@ female,������������������������       �                     �?male,30�       �                   �@      �?              @ le,10,0������������������������       �                     @ ,0,0,34�       �                 �?�@���Q��?             @ A/5. 13������������������������       �                     �? 5082,7.�       �                 ��I @      �?             @aria Br�       �                   �?@�q�q�?             @ . Vikto������������������������       �                     �?, Mr. P������������������������       �      �?              @Mrs. Cha������������������������       �                     �?,1,2,"P�       �                   @E@�J�T�?-            �Q@Marshal�       �                 �?�@�X�<ݺ?             B@ s",male������������������������       �        
             1@ mbisky)�       �                 @3�@�KM�]�?             3@ strom-S������������������������       ��q�q�?             @52,S
43�       �                   @D@      �?             0@,female������������������������       �                     ,@der (Ali�       �                     @      �?              @ ,"Kalli������������������������       �                     �? 5,,S
43������������������������       �                     �? E44,S
4������������������������       �                    �A@ 20,B96 �       �                     �?X��ʑ��?            �E@male,21�       �                 ��yC@j���� �?             A@(Emily �       �                   �A@����X�?             <@Mr. Mar�       �                 �T!@@�q�q�?             8@ Mr. Jo�       �                   �J@���!pc�?             6@1,1,2,"�       �                 `fF<@�t����?	             1@1,F.C.C�       �                 �|�?@$�q-�?             *@ 5769,9.������������������������       �                     �?76,7.77������������������������       �                     (@30434,13�       �                   @>@      �?             @ ,65306,������������������������       �                     �?,33638,8������������������������       �                     @female,�       �                 `fF<@z�G�z�?             @r",male������������������������       �                     @herine"������������������������       �                     �?thur Go������������������������       �                      @ Edwy Ar������������������������       �                     @r. Ingv������������������������       �                     @an, Mr.�       �                    ;@�<ݚ�?             "@ 1,1,"Go�       �                 ��?P@�q�q�?             @ 55,0,3,������������������������       �                      @ "Jalsev������������������������       �                     �? t, Mr. ������������������������       �                     @nyon, Mr�       �                   �:@DX�\��?3            �Q@ 459,1,2�       �                    �?��2(&�?             6@
460,0,�       �                     @     ��?             0@ 1,"Ande�       �                    2@����X�?             @ orley, ������������������������       �                     �? Arthur�       �                     �?r�q��?             @ acob Ch������������������������       �                      @Simon",m�       �                    �?      �?             @ Estansl������������������������       �                     �?bell, Mr������������������������       �                     @ Montgo�       �                   �!@�����H�?             "@ ames",m�       �                 ��Y@      �?             @ rbara",������������������������       �                     @ r",male������������������������       �                     �?0,31508������������������������       �                     @th)",fe������������������������       �                     @n S (Ma�       �                    �?Rg��J��?%            �H@ 917,D,C�       �                   @C@���|���?             &@,9.8375�       �                    �?�z�G��?             $@5,52,A1������������������������       �                     @ 1,,S
47������������������������       �                     @8,,S
479������������������������       �                     �? 8,,S
48�                           @      �?             C@2875,,S�                         @D@��}*_��?             ;@144,46.�                           �?�<ݚ�?             2@,0,2398�                       �|Y=@r�q��?	             (@ 5 3594,                       ���M@      �?              @ 34,9.58������������������������       �                     �?        ������������������������       �                     �?                                 �?ףp=
�?             $@       ������������������������       �                     @                              `f�K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                �@@�q�q�?             @       	      
                  �<@z�G�z�?             @        ������������������������       �                     �?                                �7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                  �?�q�q�?             "@                             �CdQ@      �?              @        ������������������������       �                     @                                 �?���Q��?             @        ������������������������       �                      @                              ��#[@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?"pc�
�?             &@                              ���.@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @              (                    @�^�����?R             _@                                 �? i���t�?$            �H@       ������������������������       �                     C@               !                   �?�eP*L��?             &@        ������������������������       �                     �?        "      '                   �?���Q��?             $@       #      $                    �?X�<ݚ�?             "@        ������������������������       �                      @        %      &                   :@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        )      4                   �?��n�?.            �R@        *      +                  �7@���Q��?            �A@        ������������������������       �                     (@        ,      1                ��T?@���}<S�?             7@       -      0                   @@�}�+r��?             3@        .      /                �|Y>@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             ,@        2      3                ���A@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     D@        �t�bh�h*h-K ��h/��R�(KM5KK��h]�BP       �{@     �p@     �P@     @R@      @     �K@      �?     �F@              E@      �?      @      �?                      @      @      $@      @      "@      @      @              @      @               @      @       @       @               @       @                      @              �?      N@      2@      J@      2@      J@      .@      J@      ,@     �G@      &@     �E@      $@      C@      "@      =@      "@      ;@      @      6@      @      �?      �?      �?                      �?      5@      @      &@      �?      @      �?      �?              @      �?              �?      @              @              $@      @              �?      $@      @      �?              "@      @      @      @      �?              @      @      @              @               @      @              @       @              "@              @      �?              �?      @              @      �?              �?      @              @      @      �?      @      �?      �?              �?      �?                       @      @                      �?              @       @             �w@      h@     �s@     �`@     �p@     �Z@      .@      N@      "@      ,@      @      *@      @      @              �?      @      @      @      @              �?      @       @       @       @              �?       @      �?       @                      �?      �?              �?      @              �?      �?       @              �?      �?      �?              �?      �?                      @      @      �?      �?              @      �?       @      �?              �?       @               @              @      G@              $@      @      B@       @     �@@      �?      @              @      �?              �?      >@              *@      �?      1@              "@      �?       @      �?      @      �?                      @              @      @      @              @      @              p@      G@     `m@      8@     �d@      6@     @d@      1@      W@      @     �A@      @      4@      @      4@       @      �?              3@       @      (@              @       @      �?       @      �?                       @      @                      @      .@             �L@      �?     �J@      �?      &@              E@      �?      6@              4@      �?      @      �?      0@              @             �Q@      &@      ,@      @      "@      �?      �?      �?      �?                      �?       @              @      @      @       @      �?       @      @                       @      L@      @      �?             �K@      @      6@             �@@      @      .@              2@      @      &@      �?      @              @      �?       @              @      �?              �?      @              @      @      �?      @               @      �?       @               @      �?              @      �?      @                      �?      @      @      �?              @      @              @      @       @      �?               @       @      �?       @              �?      �?      �?      �?             @Q@       @      A@       @      1@              1@       @       @      �?      .@      �?      ,@              �?      �?              �?      �?             �A@              5@      6@      ,@      4@       @      4@       @      0@      @      0@       @      .@      �?      (@      �?                      (@      �?      @      �?                      @      @      �?      @                      �?       @                      @      @              @       @      �?       @               @      �?              @              E@      =@      3@      @      *@      @      @       @              �?      @      �?       @              @      �?              �?      @               @      �?      @      �?      @                      �?      @              @              7@      :@      @      @      @      @              @      @              �?              3@      3@      $@      1@      @      ,@       @      $@      �?      �?              �?      �?              �?      "@              @      �?       @      �?                       @       @      @      �?      @              �?      �?      @      �?                      @      �?              @      @      @      @      @               @      @               @       @      �?       @                      �?      �?              "@       @      �?       @      �?                       @       @             �P@      M@      @      F@              C@      @      @      �?              @      @      @      @       @               @      @              @       @                      �?     �N@      ,@      5@      ,@              (@      5@       @      2@      �?      @      �?      @                      �?      ,@              @      �?              �?      @              D@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ$�phG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtK�huh*h-K ��h/��R�(KK���h|�B@?         .                   �3@�L*�<�?�           8�@     �F@       +                    @b�L�4��?P            �`@                                  �?�Sb(�	�?A             [@                                   �?���.�6�?             G@        ������������������������       �        
             2@                                   @ �Cc}�?             <@       ������������������������       �                     2@     @       	                    @�z�G��?             $@      �?������������������������       �                     @        
                           �?      �?             @     ?@                           �?      �?             @     @������������������������       �                     @      @������������������������       �                     �?      �?������������������������       �                      @      @                        �?�@�g�y��?#             O@        ������������������������       �                     ,@      ,@                           �?      �?             H@      �?������������������������       �                      @     �`@                            �?�LQ�1	�?             G@      *@                           �?և���X�?             <@     @                            @      �?
             8@      �?                          �2@      �?             @        ������������������������       �                      @      �?                          �'@      �?             @      @������������������������       �                     @      �?������������������������       �                     �?      G@                        ��Y @      �?             2@     @                           1@ףp=
�?             $@      *@������������������������       �      �?             @      @������������������������       �                     @      @������������������������       �                      @      8@������������������������       �                     @      @!       "                    �?�<ݚ�?             2@       @������������������������       �                      @      �?#       $                 03{3@      �?             0@        ������������������������       �                     $@        %       *                    �?�q�q�?             @     4@&       )                    �?���Q��?             @     $@'       (                    7@      �?             @        ������������������������       �                      @      3@������������������������       �                      @      @������������������������       �                     �?      �?������������������������       �                     �?      �?,       -                   -@$�q-�?             :@       @������������������������       �                      @        ������������������������       �                     8@      @/       p                    �?B�����?_           �@      @0       A                     @tHN�?q             f@     �?1       >                   @L@X'"7��?H             [@       2       3                    �?T��,��?D            @Y@      "@������������������������       �                     A@        4       =                    �?�����?-            �P@      @5       6                   �B@@4և���?             E@     �?������������������������       �                     =@        7       8                   @C@�θ�?	             *@      �?������������������������       �                     �?      @9       :                     �?r�q��?             (@      �?������������������������       �                     @       @;       <                    �?����X�?             @     �?������������������������       �                     @        ������������������������       �                      @      &@������������������������       �                     9@        ?       @                   �L@����X�?             @        ������������������������       �                      @      �?������������������������       �                     @      �?B       m                    @\X��t�?)            @Q@     �?C       l                 03�:@p�EG/��?%            �O@     @D       S                    �?d��0u��?"             N@      @E       R                    �?������?             >@     �?F       Q                 ��.@l��
I��?             ;@     @G       H                 �|Y=@X�<ݚ�?	             2@       @������������������������       �                     �?     @I       N                    �?��.k���?             1@       @J       M                    �?�<ݚ�?             "@       K       L                 X�x&@�q�q�?             @        ������������������������       �                      @       ������������������������       �                     @        ������������������������       �                     @        O       P                 �&�@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@       ������������������������       �                     @        T       k                   @B@��S���?             >@       U       f                    �?�5��?             ;@       V       ]                    �?      �?             4@       W       Z                 ��� @��
ц��?             *@       X       Y                   �9@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        [       \                    ;@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ^       _                 ���)@և���X�?             @        ������������������������       �                      @        `       e                 03�1@���Q��?             @       a       d                   �0@      �?             @       b       c                 �|�;@      �?              @        ������������������������       �                     �?       ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?       g       h                    �?؇���X�?             @        ������������������������       �                     @        i       j                 �|�:@�q�q�?             @        ������������������������       �                      @       ������������������������       �                     �?        ������������������������       �                     @       ������������������������       �                     @        n       o                 ���4@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        q       �                 ��D:@\���(\�?�             y@       r       �                    �?\2R}�?�            r@        s       ~                 �|Y=@�θV�?,            @Q@        t       }                    �?����X�?
             ,@       u       z                    �?�q�q�?             (@       v       w                   �8@�z�G��?             $@        ������������������������       �                     @        x       y                   @@      �?             @        ������������������������       �                     �?       ������������������������       �                     @       {       |                    ;@      �?              @        ������������������������       �                     �?       ������������������������       �                     �?       ������������������������       �                      @              �                 �|�=@�1�`jg�?"            �K@       �       �                    �?Du9iH��?            �E@        �       �                    �?$�q-�?
             *@.275,,S������������������������       �        	             (@v�X  ������������������������       �                     �?%��X  �       �                   `3@��S�ۿ?             >@?�X  �       �                 ���@h�����?             <@ emale,4������������������������       �                     $@female,1�       �                   @'@�X�<ݺ?
             2@Mary Hi������������������������       �$�q-�?             *@ Mr. Pet������������������������       �                     @�l�X  �       �                    �?      �?              @ :�X  ������������������������       �                     �? en, Mr.������������������������       �                     �? C�X  ������������������������       �                     (@ft, Mrs.�       �                   @4@�2�~w�?�            �k@ 7466,25�       �                 pf� @      �?             0@ ,female�       �                    �?      �?              @male,24������������������������       �                     @��X  ������������������������       �                     @ male,27������������������������       �                      @hington �       �                   �<@ =[y��?y            �i@ van Mel������������������������       �        '            @P@ �X  �       �                   �*@��X�-�?R            `a@��X  �       �                     @�#-���?@            @Z@ ckwith,�       �                   �F@r�q��?             8@U�X  �       �                   @D@���y4F�?             3@,695,5,�       �                 `fF)@r�q��?             2@E�X  ������������������������       �                     $@y)",fema�       �                 �|�=@      �?              @ ��X  ������������������������       �                      @ r. Alfr�       �                    @@r�q��?             @ r. Nede������������������������       �                     @ ��X  �       �                   @B@�q�q�?             @ (Lily ������������������������       �      �?              @1,2,"She������������������������       �                     �? ��X  ������������������������       �                     �?8958,,S
������������������������       �                     @ ,10.516�       �                 ���"@xdQ�m��?/            @T@C.A./SO�       �                 ��@ �\���?-            �S@ ?�X  ������������������������       �                     7@ ret Nor�       �                 ��L@@4և���?!             L@ ev. Juo�       �                 �|Y>@���Q��?             @ aret Ed������������������������       �                      @ ��X  ������������������������       �                     @ 90,1,1,�       �                   �@@`'�J�?            �I@�X  �       �                 ��) @`Jj��?             ?@� �0�u �       �                 @3�@h�����?             <@^�X  �       �                 �?�@��S�ۿ?             .@��X  ������������������������       �                     $@       ������������������������       �z�G�z�?             @        ������������������������       �                     *@�$�X  �       �                 �|Y=@�q�q�?             @ ��X  ������������������������       �                     �?i��X  �       �                 �|�>@      �?              @        ������������������������       �                     �?I|�X  ������������������������       �                     �?       ������������������������       �        	             4@��X  �       �                    ?@      �?              @        ������������������������       �                     �?�%�X  ������������������������       �                     �?M�X  ������������������������       �                     A@       �       �                 p�w@�/e�U��?A            �[@^�X  �       �                    �?� �W�??            �Z@q�X  �       �                    �?X�Cc�?4             U@ &�X  �       �                 @�pX@
;&����?             7@��X  �       �                    �?b�2�tk�?             2@       �       �                 �|�;@�eP*L��?             &@        ������������������������       �                      @��X  �       �                 ��2>@�q�q�?             "@ �X  ������������������������       �                      @       �       �                    C@؇���X�?             @       ������������������������       �                     @ �X  �       �                 �D D@�q�q�?             @ ��X  ������������������������       �                     �? p�X  ������������������������       �                      @        �       �                 ��`E@؇���X�?             @ 9�X  ������������������������       �                     �?        ������������������������       �                     @���X  ������������������������       �                     @ @�X  �       �                    R@�ɞ`s�?%            �N@��X  �       �                 03k:@�c�Α�?$             M@        ������������������������       �                      @        �       �                 �!fK@      �?#             L@       �       �                     �?z�G�z�?             D@       �       �                    <@��G���?            �B@ 3�X  ������������������������       �                     �? ��X  �       �                   �F@r�q��?             B@��X  �       �                    �?�E��ӭ�?             2@4�X  �       �                   `@@�n_Y�K�?
             *@        �       �                 �|Y=@r�q��?             @ l�X  ������������������������       �                     �? ��X  ������������������������       �                     @��X  ������������������������       �                     @S3�X  ������������������������       �                     @C�X  �       �                   @J@�X�<ݺ?
             2@ ��X  �       �                 `f�;@      �?              @        ������������������������       �                     �? .�X  ������������������������       �                     @        ������������������������       �                     $@��X  ������������������������       �                     @       �       �                    �?     ��?             0@       �       �                     @�n_Y�K�?	             *@       �       �                    C@�<ݚ�?             "@��X  �       �                 �|Y>@���Q��?             @       ������������������������       �                     @�.�X  ������������������������       �                      @        ������������������������       �                     @        �       �                    >@      �?             @       �       �                    ;@      �?              @ ��X  ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @8s�X  �       �                 ���[@�q�q�?             @ ��X  ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @��X  �       �                     �?�nkK�?             7@       �       �                    �?�8��8��?             (@        �       �                 ��UO@؇���X�?             @ L�X  ������������������������       �                     @        �       �                   @D@�q�q�?             @ \�X  ������������������������       �                     �?�)�X  ������������������������       �                      @        ������������������������       �                     @       ������������������������       �                     &@��X  ������������������������       �                     @       �t�b�     h�h*h-K ��h/��R�(KK�KK��h]�B�       p{@      q@     �M@     �R@     �A@     @R@      @     �E@              2@      @      9@              2@      @      @              @      @      @      �?      @              @      �?               @              @@      >@      ,@              2@      >@       @              0@      >@      (@      0@      (@      (@      @      @       @              �?      @              @      �?              "@      "@      �?      "@      �?      @              @       @                      @      @      ,@       @               @      ,@              $@       @      @       @      @       @       @       @                       @              �?              �?      8@       @               @      8@             �w@     �h@     �A@     �a@      @     �Y@      @     �X@              A@      @      P@      @     �C@              =@      @      $@      �?               @      $@              @       @      @              @       @                      9@       @      @       @                      @      >@     �C@      9@      C@      6@      C@       @      6@       @      3@       @      $@              �?       @      "@      @       @      @       @               @      @              @              �?      @      �?                      @              "@              @      ,@      0@      &@      0@      $@      $@      @      @      @       @               @      @              �?      @      �?                      @      @      @       @               @      @      �?      @      �?      �?      �?                      �?               @      �?              �?      @              @      �?       @               @      �?              @              @              @      �?              �?      @             �u@     �K@     �p@      4@      O@      @      $@      @       @      @      @      @      @              �?      @      �?                      @      �?      �?      �?                      �?       @              J@      @      D@      @      (@      �?      (@                      �?      <@       @      ;@      �?      $@              1@      �?      (@      �?      @              �?      �?      �?                      �?      (@             �i@      *@      (@      @      @      @      @                      @       @             `h@      "@     @P@             @`@      "@      X@      "@      4@      @      .@      @      .@      @      $@              @      @               @      @      �?      @               @      �?      �?      �?      �?                      �?      @              S@      @     �R@      @      7@              J@      @      @       @               @      @             �H@       @      =@       @      ;@      �?      ,@      �?      $@              @      �?      *@               @      �?      �?              �?      �?              �?      �?              4@              �?      �?              �?      �?              A@              S@     �A@      S@      ?@      K@      >@      (@      &@      @      &@      @      @               @      @      @               @      @      �?      @               @      �?              �?       @              �?      @      �?                      @      @              E@      3@      E@      0@               @      E@      ,@     �@@      @      >@      @              �?      >@      @      *@      @       @      @      �?      @      �?                      @      @              @              1@      �?      @      �?              �?      @              $@              @              "@      @       @      @      @       @      @       @      @                       @      @              �?      @      �?      �?              �?      �?                       @      �?       @      �?                       @              @      6@      �?      &@      �?      @      �?      @               @      �?              �?       @              @              &@                      @�t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJW:+LhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM)huh*h-K ��h/��R�(KM)��h|�B@J         r                    �?]@f�
�?�           8�@               a                    �?��K�"�?�            �q@              &                 `f�$@�e�U��?�            �m@      @       %                    �?��H�}�?              I@              "                    �?(���@��?            �G@                               �̌@���� �?            �D@     �?                        ���@�r����?             >@     �E@       	                 �|Y:@����X�?             @       @������������������������       �                     @        
                           �?�q�q�?             @        ������������������������       �                     �?p�X�X  ������������������������       �                      @p�X�X                             �?���}<S�?             7@�X�X  ������������������������       �        	             0@p�X�X                             4@����X�?             @ �X�X  ������������������������       �                     �?��X�X                          �&B@r�q��?             @�X                            �7@�q�q�?             @ ��X  ������������������������       �                      @P��X  ������������������������       �                     �?��X  ������������������������       �                     @P��X                            �2@���|���?             &@ ��X  ������������������������       �                     �?��X                          ��� @�z�G��?             $@��X                          @3�@r�q��?             @��X                            �8@�q�q�?             @ ��X  ������������������������       �                     �?P��X                             ;@      �?              @ ��X  ������������������������       �                     �? ��X  ������������������������       �                     �?���X  ������������������������       �                     @P��X          !                  SE"@      �?             @ ��X  ������������������������       �                      @       @������������������������       �                      @        #       $                   �3@�q�q�?             @        ������������������������       �                      @      �?������������������������       �                     @        ������������������������       �                     @      �?'       `                 �QD@X�E)9�?v            �g@       (       E                    �?�<�}���?K            @^@       )       D                    @�? Da�?(            �O@     @*       +                    �?\#r��?&            �N@      @������������������������       �                     @        ,       5                 `f�)@ �Cc}�?#             L@      @-       .                 pF%@`2U0*��?             9@       @������������������������       �                     *@      �?/       0                    +@�8��8��?             (@      @������������������������       �                     @       @1       4                    �?r�q��?             @      @2       3                 ��&@z�G�z�?             @      �?������������������������       �                     �?      �?������������������������       �                     @      4@������������������������       �                     �?      .@6       =                   �*@�חF�P�?             ?@      @7       <                   �B@X�<ݚ�?             "@       8       ;                    �?����X�?             @       9       :                    <@�q�q�?             @        ������������������������       �                      @      @������������������������       �                     @        ������������������������       �                     �?      �?������������������������       �                      @        >       ?                    �?���7�?             6@     @������������������������       �                     .@      3@@       C                    1@؇���X�?             @     �?A       B                    "@�q�q�?             @     �?������������������������       �                      @     �?������������������������       �                     �?     @������������������������       �                     @      @������������������������       �                      @     �?F       _                   �@@V�a�� �?#             M@     @G       H                    �?F�t�K��?"            �L@       @������������������������       �        	             .@     @I       J                   �9@0,Tg��?             E@       @������������������������       �                     ,@       K       T                     @��>4և�?             <@       L       M                    6@      �?             0@        ������������������������       �                      @        N       S                    :@؇���X�?
             ,@       O       P                   �8@�<ݚ�?             "@        ������������������������       �                     �?        Q       R                   �E@      �?              @       ������������������������       �                     @       ������������������������       �                      @        ������������������������       �                     @       U       ^                 �̤=@�q�q�?             (@       V       ]                 `fV6@�z�G��?             $@       W       X                 �|�;@և���X�?             @        ������������������������       �                     @        Y       Z                 03�1@      �?             @        ������������������������       �                      @        [       \                 03C3@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?       ������������������������       �        +             Q@       b       q                    @v�2t5�?            �D@       c       d                    �?      �?             A@        ������������������������       �                     @        e       f                     @�f7�z�?             =@        ������������������������       �                     @       g       h                    @�q�q�?             8@        ������������������������       �                     @        i       n                    *@p�ݯ��?
             3@       j       k                    @�8��8��?             (@        ������������������������       �                     @        l       m                    @r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        o       p                 ���4@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?       ������������������������       �                     @        s       �                 ��D:@���<��?           �z@       t       y                    $@�%�P��?�            �t@        u       v                     @"pc�
�?             &@        ������������������������       �                     @        w       x                 ��|2@����X�?             @       ������������������������       �                     @        ������������������������       �                      @       z       �                     @ E�+0+�?�            �s@        {       |                   �)@�(\����?1             T@        ������������������������       �                    �A@       }       �                 ��,@`Ӹ����?            �F@       ~                        �|�<@$�q-�?             :@        ������������������������       �                     ,@       �       �                 �|�=@r�q��?             (@        ������������������������       �                     �?,0,3,"K�       �                   �A@�C��2(�?             &@�W�X  �       �                    @@r�q��?             @ �W�X  ������������������������       �                      @ xW�X  ������������������������       �      �?             @W",femal������������������������       �                     @ . Ander������������������������       �                     3@ 2,31.27�       �                    �?��5Վ3�?�            �m@  310130�       �                    �?^������?            �A@�W�X  �       �                    �?�c�Α�?             =@tW�X  �       �                 ���@      �?             8@ 12,8.05������������������������       �                     @|W�X  �       �                   @@�q�q�?
             2@ ,S
618,�       �                   �5@X�<ݚ�?             "@ ale,26,������������������������       �                      @se",fema�       �                 �|=@և���X�?             @ e,26,0,������������������������       �                      @��W�X  ������������������������       ����Q��?             @1,0,117�       �                 �|�;@�����H�?             "@ 653,15.�       �                   �2@      �?             @ ,350029������������������������       �                     @ TW�X  ������������������������       �                     �?�:X�X  ������������������������       �                     @le,57,0,�       �                 �&�)@���Q��?             @ �W�X  ������������������������       �                      @ tcho",m������������������������       �                     @~W�X  �       �                 ��y&@�q�q�?             @ n Henry������������������������       �                      @��W�X  ������������������������       �                     @ Maeglin�       �                   @@@ ��fί�?�            `i@. Willi�       �                    �?3��e��?j            �d@1X�X  �       �                   �:@$s��O�?Z            �a@ ",femal�       �                   �2@�FVQ&�?,            �P@ ",male,�       �                   �1@      �?
             (@8W�X  �       �                   �0@�<ݚ�?             "@a (Mari�       �                 pf�@����X�?             @ ,"Thorn������������������������       �                      @ Jensen,�       �                 pFD!@���Q��?             @ �V�X  ������������������������       ��q�q�?             @Skoog, M������������������������       �                      @,3,"Foo,������������������������       �                      @ Miss. E�       �                 ���@�q�q�?             @ X�X  ������������������������       �                     �? or, Mr.�       �                 ��Y @      �?              @ ?W�X  ������������������������       �                     �?,3,"Will������������������������       �                     �?P�W�X  �       �                    �?@3����?"             K@ X�X  ������������������������       �                      @Doling,�       �                 ���@ pƵHP�?!             J@  Mr. Jo�       �                    7@z�G�z�?             @ _W�X  ������������������������       �                      @�X�X  �       �                   �8@�q�q�?             @ �U�X  ������������������������       �                     �?3.5,,S
6������������������������       �                      @ �W�X  ������������������������       �                    �G@5.5,,Q
6�       �                 ��) @��A��?.            �R@8X�X  �       �                 @3�@lGts��?$            �K@275,D48�       �                   �>@(L���?            �E@�V�X  �       �                 �|Y=@     ��?             @@ �V�X  �       �                    �?z�G�z�?             @ 5875,E5������������������������       �                     �?�W�X  ������������������������       �                     @ �W�X  �       �                 ��(@�>����?             ;@`W�X  �       �                 03�@      �?             0@ :W�X  ������������������������       �                     @993,7.77������������������������       �"pc�
�?             &@,,S
670,������������������������       �                     &@PpV�X  �       �                   �?@���!pc�?             &@ UW�X  �       �                 pff@�q�q�?             @ ,0,1,"D������������������������       �                     @3,0,2,"������������������������       �                      @ 7R�X  �       �                 �?�@z�G�z�?             @ X�X  ������������������������       �                      @ �W�X  ������������������������       ��q�q�?             @ 0,3,"Sa������������������������       �                     (@ sW�X  �       �                 ��)"@p�ݯ��?
             3@ 679,0,3�       �                 �|Y<@      �?              @ �W�X  ������������������������       �                     @PzW�X  �       �                 pf� @�q�q�?             @ �W�X  ������������������������       �                     �? ,male,2������������������������       �                      @ Anderso�       �                    �?�C��2(�?             &@ s Edwar������������������������       �                      @s Willia�       �                    (@�����H�?             "@ nW�X  �       �                   �<@z�G�z�?             @ :R�X  ������������������������       �                      @<R�X  �       �                 �|Y=@�q�q�?             @ �V�X  ������������������������       �                     �? ,S
690,������������������������       �                      @�W�X  ������������������������       �                     @:W�X  �       �                    �? 7���B�?             ;@XW�X  ������������������������       �                     6@mW�X  �       �                    �?z�G�z�?             @ �X  ������������������������       �                     �?��W�X  ������������������������       �                     @ ,male,4������������������������       �                     B@�gW�X  �                          �J@*Mp����?J            �Y@orland"�       �                 ��";@|jq��?<            �T@ +X�X  �       �                 03k:@      �?              @ 1,1,"As������������������������       �                     �?18,1,0,P�       �                 �|�?@����X�?             @ cer Vic������������������������       �                     �?0�W�X  �       �                    �?r�q��?             @  Mr. Ma������������������������       �                      @ iW�X  �       �                   �C@      �?             @ ry Samu������������������������       �                     �? 1,2,"Ke�       �                    H@�q�q�?             @,S
708,������������������������       �      �?              @ �W�X  ������������������������       �                     �?113781,1�       �                   �;@L�qA��?5            �R@ am Geor�       �                    6@l��[B��?             =@�W�X  �       �                    �?�����?             3@�W�X  ������������������������       �                     "@24,S
71�       �                    @���Q��?             $@ 6,S
714������������������������       �                     @FX�X  �       �                    @�q�q�?             @,0,3,"S�       �                    @���Q��?             @ 8124,7.������������������������       �                      @��W�X  ������������������������       �                     @ ia ""Wi������������������������       �                     �?��W�X  �       �                    �?ףp=
�?             $@bW�X  ������������������������       �                     "@Annie Je������������������������       �                     �?, Mr. Sv�                           �?���j��?!             G@5X�X  �                         �I@P����?             C@ Mr. He�                          �?<ݚ)�?             B@SW�X  �                         �H@����X�?            �A@ic, Mr.                       p�w@     ��?             @@ Peter                          �?������?             >@                             `f�B@�GN�z�?             6@                               �A@�eP*L��?	             &@             	                   �?�q�q�?             "@                              �|�=@�q�q�?             @        ������������������������       �                     �?                                �A@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        
                        �>@r�q��?             @                               @=@�q�q�?             @        ������������������������       �                     �?                              �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     &@                                 �?      �?              @                             `ށK@և���X�?             @        ������������������������       �                      @                                �G@���Q��?             @                                @C@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        !      (                   �?�}�+r��?             3@       "      #                   �?$�q-�?	             *@        ������������������������       �                     @        $      '                 )?@r�q��?             @        %      &                  �Q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h*h-K ��h/��R�(KM)KK��h]�B�       z@     `r@      O@     @k@      C@      i@      2@      @@      .@      @@      &@      >@      @      :@       @      @              @       @      �?              �?       @               @      5@              0@       @      @      �?              �?      @      �?       @               @      �?                      @      @      @              �?      @      @      @      �?       @      �?      �?              �?      �?              �?      �?              @               @       @               @       @              @       @               @      @              @              4@      e@      4@     @Y@       @     �K@      @     �K@              @      @      I@      �?      8@              *@      �?      &@              @      �?      @      �?      @      �?                      @              �?      @      :@      @      @       @      @       @      @       @                      @              �?       @              �?      5@              .@      �?      @      �?       @               @      �?                      @       @              (@      G@      &@      G@              .@      &@      ?@              ,@      &@      1@      @      (@       @               @      (@       @      @              �?       @      @              @       @                      @      @      @      @      @      @      @      @              �?      @               @      �?      �?      �?                      �?      @                       @      �?                      Q@      8@      1@      1@      1@              @      1@      (@              @      1@      @      @              (@      @      &@      �?      @              @      �?              �?      @              �?      @              @      �?              @             0v@      S@      r@     �D@       @      "@              @       @      @              @       @             �q@      @@     �S@       @     �A@             �E@       @      8@       @      ,@              $@       @              �?      $@      �?      @      �?       @              @      �?      @              3@              j@      >@      7@      (@      5@       @      2@      @      @              (@      @      @      @               @      @      @       @               @      @       @      �?      @      �?      @                      �?      @              @       @               @      @               @      @       @                      @      g@      2@     �b@      2@     �^@      1@      O@      @      "@      @      @       @      @       @       @              @       @      �?       @       @               @               @      �?      �?              �?      �?              �?      �?             �J@      �?       @             �I@      �?      @      �?       @               @      �?              �?       @             �G@             �N@      *@     �H@      @     �B@      @      =@      @      @      �?              �?      @              9@       @      ,@       @      @              "@       @      &@               @      @      @       @      @                       @      @      �?       @               @      �?      (@              (@      @       @      @              @       @      �?              �?       @              $@      �?       @               @      �?      @      �?       @               @      �?              �?       @              @              :@      �?      6@              @      �?              �?      @              B@             �P@     �A@     �H@      A@       @      @              �?       @      @      �?              �?      @               @      �?      @              �?      �?       @      �?      �?              �?     �G@      <@      ,@      .@      *@      @      "@              @      @              @      @       @      @       @               @      @              �?              �?      "@              "@      �?             �@@      *@      9@      *@      9@      &@      9@      $@      6@      $@      6@       @      1@      @      @      @      @      @      �?       @              �?      �?      �?      �?                      �?      @      �?       @      �?      �?              �?      �?      �?                      �?      @                       @      &@              @      @      @      @       @               @      @       @      �?              �?       @                       @      �?                       @      @                      �?               @       @              2@      �?      (@      �?      @              @      �?      �?      �?      �?                      �?      @              @        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJF<KdhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtM'huh*h-K ��h/��R�(KM'��h|�B�I                             @	dm#��?�           8�@                                   @     ��?              H@                               �-]@(;L]n�?             >@     (@������������������������       �                     <@       @                        �(\�?      �?              @ will be������������������������       �                     �? turns
 ������������������������       �                     �?essions        	                    �?�<ݚ�?
             2@ ch valu������������������������       �                     $@      $@
                        ��T?@      �?              @        ������������������������       �                      @       @                           @�q�q�?             @    �a@������������������������       �                     @      P@������������������������       �                      @               "                  @L@^ɼ���?�           ��@     @       W                    �?@\L5�T�?�           ؃@               4                     @l��TO��?H            @_@     �?                           �?�M���?(             Q@     �`@                        03�=@�X�<ݺ?             B@      *@                            �?      �?              @      @������������������������       �                      @      �?������������������������       �                     @        ������������������������       �                     <@      �?       )                 �D�G@     ��?             @@     @                          �;@��.k���?             1@      �?������������������������       �                     �?      G@       (                     �?     ��?
             0@     @       '                    �?��
ц��?             *@     *@       &                    C@�q�q�?             (@     @       %                   �A@�eP*L��?             &@     @       $                 ��2>@���Q��?             $@     8@        #                 �ܵ<@      �?              @     @!       "                 X�,@@      �?             @       @������������������������       �                      @      �?������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @     4@������������������������       �                     �?     $@������������������������       �                     �?        ������������������������       �                     �?      3@������������������������       �                     @      @*       +                  �}S@������?
             .@      �?������������������������       �                     @      �?,       3                    �?      �?              @      @-       2                    �?�q�q�?             @       .       1                    �?      �?             @     @/       0                   �=@�q�q�?             @      @������������������������       �                     �?     �?������������������������       �                      @       ������������������������       �                     �?      "@������������������������       �                      @        ������������������������       �                      @      @5       N                    �?�MWl��?             �L@     �?6       9                    �?:	��ʵ�?            �F@        7       8                 `�@1@      �?              @     �?������������������������       �                     @      @������������������������       �                      @      �?:       G                 �|Y=@�MI8d�?            �B@       @;       @                 ���@X�Cc�?             ,@      �?<       =                    5@���Q��?             @        ������������������������       �                     �?      &@>       ?                   �7@      �?             @        ������������������������       �                     @        ������������������������       �                     �?      �?A       F                   �<@�<ݚ�?             "@     �?B       C                   �8@      �?              @      �?������������������������       �                     @     @D       E                   @;@�q�q�?             @      @������������������������       �                     �?     �?������������������������       �                      @     @������������������������       �                     �?       @H       I                 ���@�nkK�?             7@      @������������������������       �                     @       @J       M                 �|�=@      �?             0@       K       L                   @@�C��2(�?             &@       ������������������������       �؇���X�?             @        ������������������������       �                     @        ������������������������       �                     @       O       V                 ���.@�q�q�?             (@       P       U                    �?      �?              @       Q       R                    �?r�q��?             @        ������������������������       �                     @       S       T                 �&�)@      �?              @        ������������������������       �                     �?       ������������������������       �                     �?       ������������������������       �                      @       ������������������������       �                     @        X                       0�^I@Gq����?F           �@       Y       �                     @�"��c��?           P|@        Z       �                    �?z�7�Z�?\            @b@       [       t                 �|Y=@$��fF?�?L            @_@        \       a                    &@H�z�G�?             D@        ]       ^                    �?X�Cc�?             ,@        ������������������������       �                     @        _       `                   �7@����X�?             @        ������������������������       ��q�q�?             @       ������������������������       �                     @       b       k                   �;@�	j*D�?             :@       c       f                    �?�t����?             1@        d       e                    7@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?       g       h                    :@��S�ۿ?             .@       ������������������������       �        	             (@        i       j                     �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        l       m                    �?�q�q�?             "@        ������������������������       �                     @        n       s                 `f�D@���Q��?             @       o       p                 `fF<@�q�q�?             @        ������������������������       �                     �?        q       r                   �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?       ������������������������       �                      @        u       �                   �*@ܻ�yX7�?1            @U@        v       }                   �>@��p\�?            �D@        w       x                    �?�r����?
             .@        ������������������������       �                     �?        y       |                 �|�=@@4և���?	             ,@       z       {                    @�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?       ������������������������       �                     @       ~                           �? ��WV�?             :@        ������������������������       �                     �?       ������������������������       �                     9@        �       �                   �2@���|���?             F@ ,0,3,"K������������������������       �                     @�W�X  �       �                   @J@�z�G��?             D@�W�X  �       �                    �?�q�q�?             B@xW�X  �       �                    �?`�Q��?             9@ ",femal������������������������       �                      @ . Ander�       �                     �?��+7��?             7@2,31.27�       �                   �>@�z�G��?             4@ 310130�       �                 ��<:@�eP*L��?             &@ �W�X  ������������������������       �                      @tW�X  �       �                 X��B@�q�q�?             "@ 12,8.05������������������������       �                      @|W�X  �       �                    H@և���X�?             @,S
618,������������������������       �      �?             @ ale,26,������������������������       �                     �?se",fema������������������������       �                     "@ e,26,0,������������������������       �                     @��W�X  �       �                    �?���|���?             &@ 1,0,117�       �                   �E@�q�q�?             @653,15.������������������������       �                     @ ,350029������������������������       �                      @ TW�X  ������������������������       �                     @�:X�X  ������������������������       �                     @le,57,0,�       �                    *@���N8�?             5@ �W�X  ������������������������       �                      @ tcho",m�       �                    �?�S����?             3@~W�X  ������������������������       �                     0@ n Henry������������������������       �                     @��W�X  �       �                    �?4����?�            0s@ Maeglin�       �                    �?      �?             L@ . Willi�       �                    @���B���?             :@1X�X  �       �                    �?���}<S�?             7@",femal�       �                 �|�9@      �?	             0@ ",male,������������������������       �                     @8W�X  �       �                  ��@z�G�z�?             $@ a (Mari������������������������       �                      @ ,"Thorn������������������������       �                      @ Jensen,������������������������       �                     @ �V�X  ������������������������       �                     @Skoog, M������������������������       �                     >@,3,"Foo,�       �                    �?���w;�?�            `o@ Miss. E�       �                    �?�G�5��?)            @Q@X�X  �       �                 ���1@b�2�tk�?             B@or, Mr.�       �                 �|�<@��S���?             >@?W�X  �       �                 pf�@�q�q�?             2@ 3,"Will������������������������       �                     @P�W�X  �       �                   �2@z�G�z�?	             .@ X�X  ������������������������       �                     @Doling,�       �                    �?      �?             (@ Mr. Jo�       �                   �@�<ݚ�?             "@ _W�X  �       �                 �&B@�q�q�?             @X�X  �       �                   �7@      �?              @ �U�X  ������������������������       �                     �?3.5,,S
6������������������������       �                     �? �W�X  ������������������������       �                     �?5.5,,Q
6������������������������       �                     @8X�X  �       �                 �!@�q�q�?             @ 275,D48������������������������       �                     �?�V�X  ������������������������       �                      @ �V�X  �       �                    �?�q�q�?	             (@ 5875,E5�       �                   &@      �?             @�W�X  ������������������������       �                     @ �W�X  ������������������������       �                     �?`W�X  �       �                 ��Y.@      �?              @ :W�X  ������������������������       �                     �?993,7.77������������������������       �                     @,,S
670,������������������������       �                     @PpV�X  �       �                    :@�C��2(�?            �@@UW�X  �       �                   �6@@�0�!��?
             1@,0,1,"D�       �                   �0@��S�ۿ?	             .@3,0,2,"������������������������       �                     "@ 7R�X  �       �                    3@r�q��?             @ X�X  ������������������������       �                     �? �W�X  ������������������������       �                     @ 0,3,"Sa������������������������       �                      @ sW�X  ������������������������       �                     0@ 679,0,3�       �                 �?�@|)����?z            �f@ �W�X  �       �                    ?@@�)�n�?9            @U@zW�X  �       �                    �?�\=lf�?-            �P@�W�X  �       �                 ���@ ������?)            �O@ ,male,2�       �                   �8@�����H�?             "@ Anderso�       �                   �4@z�G�z�?             @ s Edwar������������������������       �                     �?s Willia�       �                 �&b@      �?             @ nW�X  ������������������������       �                     @ :R�X  ������������������������       �                     �?<R�X  ������������������������       �                     @ �V�X  ������������������������       �        #             K@ ,S
690,������������������������       �                     @�W�X  �       �                 �&B@�����H�?             2@:W�X  ������������������������       �                     (@XW�X  �       �                   �A@�q�q�?             @ mW�X  �       �                   �@      �?             @ �X  ������������������������       �                      @��W�X  ������������������������       �                      @ ,male,4������������������������       �                      @�gW�X  �                          �?�*v��?A            @X@orland"�       �                 @3�@ ��~���?<            �V@ +X�X  �       �                    �?X�Cc�?             ,@1,1,"As�       �                   �A@�	j*D�?             *@8,1,0,P�       �                   �:@"pc�
�?             &@ cer Vic������������������������       �                     @0�W�X  ������������������������       ����Q��?             @  Mr. Ma������������������������       �                      @ iW�X  ������������������������       �                     �? ry Samu�       �                    )@�KM�]�?4             S@ 1,2,"Ke������������������������       �                     �?,S
708,�                          ?@���Lͩ�?3            �R@�W�X  �                       �|�=@H�ՠ&��?$             K@13781,1�                          �?���C��?#            �J@am Geor�                          �?�t����?!            �I@�W�X  �                       @3�!@(L���?            �E@�W�X  �       �                 �|Y<@@�0�!��?             A@24,S
71�       �                 pf� @      �?             0@6,S
714�       �                 0S5 @"pc�
�?	             &@FX�X  �       �                   �3@�<ݚ�?             "@ ,0,3,"S�       �                   �1@      �?             @ 8124,7.������������������������       �                     �?��W�X  ������������������������       ��q�q�?             @ ia ""Wi������������������������       �                     @��W�X  ������������������������       �                      @bW�X  �       �                    8@���Q��?             @nnie Je������������������������       �                     @, Mr. Sv������������������������       �                      @5X�X  �       �                 ��) @�����H�?
             2@ Mr. He������������������������       �                     .@SW�X  �                        pf� @�q�q�?             @ ic, Mr.������������������������       �                      @ Peter ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     5@        ������������������������       �                     @                                  @�q�q�?*            �L@       	      
                   �?���3�E�?%             J@       ������������������������       �                     @@                                 �?      �?             4@                                 �?�E��ӭ�?             2@                               �E@     ��?             0@                              x#J@�n_Y�K�?             *@        ������������������������       �                     @                                 �?      �?             $@        ������������������������       �                     �?                              `�iJ@X�<ݚ�?             "@        ������������������������       �                     @                              `f�N@�q�q�?             @                                7@      �?             @        ������������������������       �                     �?                                 A@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @              !                   �?z�G�z�?             @                                  ;@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        #      &                   �?h�����?             <@        $      %                  pE@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     :@        �t�bh�h*h-K ��h/��R�(KM'KK��h]�Bp       0}@     �n@      .@     �@@      �?      =@              <@      �?      �?              �?      �?              ,@      @      $@              @      @       @               @      @              @       @             @|@     `j@     �z@     @j@     �M@     �P@      .@     �J@       @      A@       @      @       @                      @              <@      *@      3@      "@       @              �?      "@      @      @      @      @      @      @      @      @      @       @      @       @       @       @                       @              @       @              �?                      �?      �?              @              @      &@              @      @      @      @       @       @       @      �?       @      �?                       @      �?               @                       @      F@      *@     �B@       @      @       @      @                       @      ?@      @      "@      @       @      @      �?              �?      @              @      �?              @       @      @      �?      @               @      �?              �?       @                      �?      6@      �?      @              .@      �?      $@      �?      @      �?      @              @              @      @      @      �?      @      �?      @              �?      �?              �?      �?               @                      @     �v@      b@     �u@     �Z@     �W@      J@     @V@      B@      7@      1@      @      "@              @      @       @      �?       @      @              2@       @      .@       @      �?      �?              �?      �?              ,@      �?      (@               @      �?              �?       @              @      @              @      @       @      �?       @              �?      �?      �?              �?      �?               @             �P@      3@      C@      @      *@       @              �?      *@      �?      $@      �?      $@                      �?      @              9@      �?              �?      9@              <@      0@              @      <@      (@      8@      (@      1@       @               @      1@      @      ,@      @      @      @       @              @      @               @      @      @      @      @              �?      "@              @              @      @       @      @              @       @              @              @              @      0@       @              @      0@              0@      @             �o@      K@     �A@      5@      @      5@       @      5@       @      ,@              @       @       @       @                       @              @      @              >@             @k@     �@@      J@      1@      6@      ,@      0@      ,@      (@      @              @      (@      @      @              "@      @      @       @      �?       @      �?      �?              �?      �?                      �?      @               @      �?              �?       @              @       @      @      �?      @                      �?      �?      @      �?                      @      @              >@      @      ,@      @      ,@      �?      "@              @      �?              �?      @                       @      0@             �d@      0@     �T@      @     �P@      �?      O@      �?       @      �?      @      �?      �?              @      �?      @                      �?      @              K@              @              0@       @      (@              @       @       @       @               @       @               @              U@      *@     @S@      *@      "@      @      "@      @      "@       @      @              @       @               @              �?      Q@       @              �?      Q@      @     �G@      @     �G@      @     �F@      @     �B@      @      <@      @      (@      @      "@       @      @       @       @       @      �?              �?       @      @               @              @       @      @                       @      0@       @      .@              �?       @               @      �?              "@               @               @                      �?      5@              @              3@      C@      .@     �B@              @@      .@      @      *@      @      &@      @       @      @      @              @      @      �?              @      @              @      @       @       @       @      �?              �?       @               @      �?               @              @               @               @              @      �?      �?      �?              �?      �?              @              ;@      �?      �?      �?      �?                      �?      :@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJؽ�hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�C         P                     �?e�L��?�           8�@    X         3                    �?�G�z�?f             d@     @                           �?���r
��?A            @X@ pñX                             �?�D����?             E@ f e s                           @H@p�ݯ��?             C@     @                        �|�;@�������?             >@       @������������������������       �                     &@      ;@       	                    �?p�ݯ��?             3@      @������������������������       �                     $@`�zO�  
                          �A@�<ݚ�?             "@�zO�                          X�,@@����X�?             @�zO�                          ��2>@r�q��?             @ �zO�  ������������������������       �                     �?(�zO�  ������������������������       �                     @�zO�  ������������������������       �                     �?0g�X  ������������������������       �                      @wkO�                          ��Z@      �?              @     �?������������������������       �                     @     �`@������������������������       �                     �?      *@                        �\@      �?             @      @������������������������       �                     �?      �?������������������������       �                     @               *                 0�_J@N{�T6�?$            �K@     �?                           �?��.k���?             A@      @������������������������       �                     @      �?                        �|�<@���Q��?             >@      G@������������������������       �                     @     @       )                    R@�q�q�?             ;@     *@       (                    L@�	j*D�?             :@     @       '                   �>@���Q��?             4@     @                         �̌*@�q�q�?             (@      8@������������������������       �                      @     @!       "                   �C@z�G�z�?             $@      (@������������������������       �                     @      @#       &                 `f�;@�q�q�?             @      @$       %                    H@z�G�z�?             @       ������������������������       �      �?             @      @������������������������       �                     �?      0@������������������������       �                     �?        ������������������������       �                      @      5@������������������������       �                     @        ������������������������       �                     �?        +       0                 03c@؇���X�?             5@     ,@,       -                    �?�IєX�?	             1@       ������������������������       �                     .@      �?.       /                    =@      �?              @        ������������������������       �                     �?       @������������������������       �                     �?      @1       2                 ���f@      �?             @      @������������������������       �                      @      �?������������������������       �                      @        4       O                   �P@�<ݚ�?%            �O@     �?5       @                 ��Q@���*�?$             N@      �?6       7                    �?�q�q�?             2@        ������������������������       �                     @       @8       ?                    F@�eP*L��?             &@       9       :                    �?r�q��?             @      @������������������������       �                      @       @;       >                   @B@      �?             @     @<       =                   @K@�q�q�?             @      @������������������������       �                     �?       @������������������������       �                      @        ������������������������       �                     �?       @������������������������       �                     @       @A       H                    �?���H��?             E@       B       G                    �?`Jj��?             ?@     C@C       D                    �?$�q-�?             :@     @������������������������       �        
             2@      @E       F                 ���^@      �?              @      @������������������������       �                     @       @������������������������       �                      @        ������������������������       �                     @      �?I       L                    �?���!pc�?             &@     �?J       K                 �U�X@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        M       N                 ��f`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        Q       �                    �?�w�+`�?]           8�@       R       �                 Ь�#@�;�T<:�?           �z@       S       T                 ���@D�a�ў�?�            �p@        ������������������������       �                     <@        U       V                 ��@�.�PI�?�            �m@        ������������������������       �                     @        W       X                    /@P�z�?�            `m@        ������������������������       �                      @        Y       p                    �?F�|���?�             m@        Z       [                    �?Dc}h��?&             L@        ������������������������       �        	             *@        \       i                    �?�ʈD��?            �E@       ]       h                 �� @�LQ�1	�?             7@       ^       a                 ���@؇���X�?             5@        _       `                 �|�9@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        b       g                 �|Y=@r�q��?	             (@        c       d                   @8@�q�q�?             @        ������������������������       �                     �?        e       f                   @@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                      @        j       k                 ���@P���Q�?             4@        ������������������������       �                     @        l       o                 X�I@      �?             0@       m       n                 ��(@��S�ۿ?             .@       ������������������������       �$�q-�?             *@        ������������������������       �                      @        ������������������������       �                     �?        q       v                    �?$���?f             f@        r       u                   �@
;&����?             7@        s       t                   �A@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                     &@        w       �                 �?�@�C��2(�?Z            @c@       x       y                 �|�<@����D��?5            @W@       ������������������������       �                     J@        z       �                   @@@������?            �D@       {       �                   �@�8��8��?             8@        |       �                 �&B@����X�?             @       }       ~                 ��@r�q��?             @        ������������������������       �                     @               �                 �|Y>@�q�q�?             @       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             1@        ������������������������       �                     1@        �       �                   �4@`��:�?%            �N@        �       �                   �0@�q�q�?
             .@        ������������������������       ����Q��?             @        �       �                 @3�@�z�G��?             $@        ������������������������       �                      @        �       �                 ��Y @      �?              @        �       �                   �2@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 @3�@*
;&���?             G@        �       �                   �A@      �?              @        ������������������������       �      �?             @        ������������������������       �      �?              @        �       �                    �?�˹�m��?             C@       �       �                 �|Y=@�8��8��?             B@        ������������������������       �                     "@        �       �                 �|Y?@�����H�?             ;@       �       �                 ��) @r�q��?	             2@       ������������������������       �                     &@        �       �                 pf� @և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                      @        �       �                   �F@v�_���?e            �c@       �       �                   P,@�S��<�?Y            �a@        �       �                    �?      �?$             N@        �       �                     @ 7���B�?             ;@       ������������������������       �                     4@        �       �                    �?؇���X�?             @       �       �                 �[$@r�q��?             @        ������������������������       �                     @        �       �                 ��&@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                 �%@<���D�?            �@@        ������������������������       �                     @        �       �                     @8�Z$���?             :@       �       �                 �|�<@�8��8��?             8@       ������������������������       �                     &@        �       �                 �|�=@8�Z$���?             *@        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                      @        �       �                 pf�/@d�� z�?5            @T@        �       �                    1@      �?             0@        �       �                   �-@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             ,@        �       �                     @�4��?)            @P@       �       �                    �?؀�:M�?            �B@        �       �                    �?      �?
             0@        ������������������������       �                     @        �       �                    �?z�G�z�?             $@        ������������������������       �                     @        �       �                   �;@����X�?             @        ������������������������       �                     �?        �       �                   �E@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@        �       �                 ���1@����X�?             <@        �       �                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                    �?R���Q�?             4@        �       �                   �2@      �?              @        ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                      @        �       �                 �|�;@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        �       �                   �.@�IєX�?             1@       ������������������������       �        	             ,@        �       �                    5@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     @X9����?U            �_@        �       �                   �6@�������?             A@        ������������������������       �        
             .@        �       �                 ��J@�\��N��?             3@       �       �                    @���Q��?             .@       �       �                    �?X�Cc�?             ,@        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?R�(��?=            @W@        �       �                 X��B@���y4F�?             3@       �       �                    @r�q��?             2@       �       �                    �?d}h���?             ,@       �       �                    3@r�q��?	             (@       �       �                    &@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                 �|Y=@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �                       �̼6@^��4m�?0            �R@        �                       �̌5@�'�=z��?            �@@       �       �                   �*@*;L]n�?             >@        �       �                    (@�z�G��?             $@       ������������������������       �                     @        �       �                 xFT$@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�z�G��?             4@       �       �                     @8�Z$���?	             *@       �       �                    )@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @        �       �                 @33/@և���X�?             @        ������������������������       �                     �?        �                           �?�q�q�?             @        ������������������������       �                     @                                 +@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @              
                   �?��p\�?            �D@              	                  @C@�t����?
             1@                                �B@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@                              ��p@@ �q�q�?             8@                              ��T?@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �        
             *@        �t�b��     h�h*h-K ��h/��R�(KMKK��h]�B�       �{@     �p@      J@      [@      C@     �M@      1@      9@      ,@      8@      @      7@              &@      @      (@              $@      @       @      @       @      @      �?              �?      @                      �?       @              @      �?      @                      �?      @      �?              �?      @              5@      A@      2@      0@              @      2@      (@              @      2@      "@      2@       @      (@       @      @       @       @               @       @              @       @      @      �?      @      �?      @              �?      �?               @              @                      �?      @      2@      �?      0@              .@      �?      �?              �?      �?               @       @       @                       @      ,@     �H@      &@     �H@      @      (@              @      @      @      �?      @               @      �?      @      �?       @      �?                       @              �?      @              @     �B@       @      =@       @      8@              2@       @      @              @       @                      @      @       @      �?      @              @      �?               @       @       @                       @      @             px@      d@     0t@     @Y@     `k@     �G@      <@             �g@     �G@              @     �g@      F@               @     �g@      E@     �C@      1@              *@     �C@      @      4@      @      2@      @       @      �?              �?       @              $@       @      �?       @              �?      �?      �?      �?                      �?      "@               @              3@      �?      @              .@      �?      ,@      �?      (@      �?       @              �?              c@      9@      (@      &@      �?      &@              &@      �?              &@             �a@      ,@     �V@       @      J@             �C@       @      6@       @      @       @      @      �?      @               @      �?      �?      �?      �?                      �?      1@              1@             �H@      (@      $@      @      @       @      @      @               @      @      �?      @      �?              �?      @              @             �C@      @      @      @      @      @      �?      �?     �A@      @     �@@      @      "@              8@      @      .@      @      &@              @      @              @      @              "@               @              Z@      K@      V@     �J@      >@      >@      �?      :@              4@      �?      @      �?      @              @      �?       @      �?                       @              �?      =@      @      @              6@      @      6@       @      &@              &@       @               @      &@                       @      M@      7@      .@      �?      �?      �?      �?                      �?      ,@             �E@      6@      7@      ,@       @      ,@              @       @       @              @       @      @      �?              �?      @              @      �?              5@              4@       @      @      @              @      @              1@      @      @      @      @               @      @               @       @      �?              �?       @              (@              0@      �?      ,@               @      �?              �?       @              Q@     �M@      "@      9@              .@      "@      $@      "@      @      "@      @              @      "@                      �?              @     �M@      A@      @      .@      @      .@      @      &@       @      $@       @      @              @       @                      @      �?      �?              �?      �?                      @      �?             �K@      3@      1@      0@      1@      *@      @      @              @      @       @      @                       @      ,@      @      &@       @      "@       @               @      "@               @              @      @      �?               @      @              @       @      �?              �?       @                      @      C@      @      .@       @      @       @      @                       @      "@              7@      �?      $@      �?      $@                      �?      *@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJX��vhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B@A         d                    �?e�L��?�           8�@  X         _                    @<�T]���?�            �o@              \                    @Q��"�?�            `m@      @       G                 �|�=@��^���?�             m@     @                           !@ܱ#_��?\            `b@        ������������������������       �                     ,@                                   '@���c�?T            �`@      "@������������������������       �                     @      �?	                            @:�����?R            �_@       @
                           �?���J��?"            �I@     @Y@������������������������       �                     4@      I@                           �?�g�y��?             ?@     @                           9@P���Q�?             4@      @                           �?      �?             @     @                          �'@      �?              @      �?������������������������       �                     �?      @������������������������       �                     �?      @������������������������       �                      @        ������������������������       �                     0@     �[@������������������������       �                     &@      2@       :                    �?���=A�?0             S@     @       %                 @� @     ��?)             P@     �?                          �6@��s����?             E@      ,@������������������������       �        
             4@      @                          �9@���|���?             6@                                pf�@      �?             @        ������������������������       �                     �?        ������������������������       �                     @      6@                           ;@�E��ӭ�?             2@      .@������������������������       �                      @               $                    �?     ��?             0@               #                 ���@d}h���?	             ,@      @!       "                 �Y�@���Q��?             @      (@������������������������       �                      @      @������������������������       �                     @      @������������������������       �                     "@       ������������������������       �                      @      @&       1                    �?8�A�0��?             6@      0@'       (                   �,@      �?             (@        ������������������������       �                      @      5@)       0                    �?�z�G��?             $@       *       /                  S�-@�q�q�?             "@       +       .                 �|Y6@���Q��?             @     ,@,       -                   �-@�q�q�?             @        ������������������������       �                     �?      �?������������������������       �                      @        ������������������������       �                      @       @������������������������       �                     @      @������������������������       �                     �?      @2       9                 �|�:@���Q��?	             $@     �?3       8                    �?؇���X�?             @       4       5                  �#@      �?             @      �?������������������������       �                      @      �?6       7                 �[$@      �?              @        ������������������������       �                     �?       @������������������������       �                     �?       ������������������������       �                     @      @������������������������       �                     @       @;       @                   �6@�q�q�?             (@      @<       ?                   �3@z�G�z�?             @     @=       >                    �?      �?             @       @������������������������       �                     @        ������������������������       �                     �?       @������������������������       �                     �?       @A       B                 �|�:@և���X�?             @        ������������������������       �                      @        C       D                    �?z�G�z�?             @        ������������������������       �                      @        E       F                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        H       W                    �?�̨�`<�?8            @U@       I       J                   @B@؇���X�?%             L@       ������������������������       �                     ;@        K       V                 83'E@�c�Α�?             =@       L       O                     �?      �?	             0@        M       N                    �?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        P       U                   �+@�<ݚ�?             "@       Q       T                     @�q�q�?             @       R       S                    D@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     *@        X       Y                     @XB���?             =@       ������������������������       �                     7@        Z       [                    C@r�q��?             @        ������������������������       �                     @        ������������������������       �                     �?        ]       ^                 ��T?@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        `       a                      @�t����?             1@        ������������������������       �                     @        b       c                 �|Y?@$�q-�?
             *@       ������������������������       �        	             (@        ������������������������       �                     �?        e       �                 ��K.@�#2����?"           �|@       f       w                    �?�]l*7��?�            0r@        g       h                   �6@>���Rp�?             M@        ������������������������       �                     "@        i       n                 �|Y=@ i���t�?            �H@        j       m                    �?      �?             (@       k       l                   �<@�q�q�?             "@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        o       p                 ���@@-�_ .�?            �B@        ������������������������       �                     .@        q       r                     @�C��2(�?             6@        ������������������������       �                     @        s       v                 �|�=@�����H�?	             2@       t       u                   @@"pc�
�?             &@       ������������������������       �����X�?             @        ������������������������       �                     @        ������������������������       �                     @        x       �                    �?`�q��־?�             m@       y       �                 ���"@ �Cc��?�             l@       z       �                 ��@�1��?o            �e@        {       |                     @��v$���?*            �N@        ������������������������       �                     $@        }       �                 ���@���J��?#            �I@        ~                        ���@�IєX�?
             1@       ������������������������       �        	             0@        ������������������������       �                     �?        ������������������������       �                     A@01310,7�       �                    �?�h����?E             \@5,,Q
36�       �                   �3@ ѯ��?B            �Z@ ,7.25,,�       �                   �1@��2(&�?             6@ n)",fem������������������������       �                     &@ oura Bo�       �                 �?�@���!pc�?             &@ Annie",������������������������       �                     @ Pauline�       �                 ��Y @���Q��?             @George �       �                   �2@      �?             @ d, Mr. ������������������������       �                      @ an, Mr.������������������������       �      �?              @ghini, M������������������������       �                     �?son, Mis�       �                 �|Y=@@�)�n�?6            @U@ yer, Mr������������������������       �                    �B@ 8,,C
37�       �                   @@@      �?             H@077,7.2�       �                    ?@�#-���?            �A@03,211.�       �                 �|�=@@4և���?             <@0125,,C�       �                  sW@HP�s��?             9@ ,7.775,������������������������       �      �?             @7,227.52������������������������       �                     5@ ,2653,1������������������������       �                     @ 2. 310�       �                 P�@؇���X�?             @ ary Ali������������������������       �                     �?ky, Mr.������������������������       �                     @ harles ������������������������       �                     *@  Master������������������������       �                     @ss, Miss�       �                   @B@�t����?$            �I@atthew"�       �                   �@@R���Q�?             D@a",fema�       �                     @�ݜ�?            �C@st",mal�       �                    5@���7�?             6@ Olof",m�       �                   �2@z�G�z�?             @ n Birge������������������������       �                      @ rjorie"������������������������       ��q�q�?             @ s. Hjal������������������������       �                     1@ .7,G6,S�       �                 `�X#@������?             1@,S
397,�       �                   �<@�	j*D�?             *@ 398,0,2������������������������       �                     @ 2,"Pain�       �                 �|Y=@X�<ݚ�?             "@ Mrs. Wi������������������������       �                      @ ,"Niska�       �                 �|�=@����X�?             @ ,0,3,"A������������������������       �                     @ la, Mis�       �                   �?@      �?             @ ainen, ������������������������       �                      @ 405,0,3������������������������       �                      @ 
406,0,������������������������       �                     @ idegren������������������������       �                     �? 1,2,"Ri������������������������       �                     &@09,0,3,�       �                    �?�<ݚ�?             "@ 775,,S
������������������������       �                      @ 411,0,3�       �                    �?����X�?             @"Hart, �       �                     @���Q��?             @ iss. Da������������������������       �                      @Mr. Alf������������������������       �                     @ Johan J������������������������       �                      @ek, Mrs�       �                   �A@      �?l             e@S
417,1�       �                   @A@�Sb(�	�?D             [@le,34,1�       �                 `�/@�Y|���?A            �Y@ female,������������������������       �                     @male,30�       �                    @�D��??            �X@le,10,0�       �                    �?^H���+�?3            �R@,0,0,34�       �                    �?�Gi����?            �B@A/5. 13�       �                    �?���|���?            �@@ 5082,7.�       �                      @�q�q�?             "@aria Br�       �                 �|Y<@����X�?             @ . Vikto�       �                    9@�q�q�?             @ , Mr. P������������������������       �                     �?Mrs. Cha������������������������       �                      @,1,2,"P������������������������       �                     @Marshal�       �                   �2@      �?              @ s",male������������������������       �                     �? mbisky)������������������������       �                     �? strom-S�       �                   �?@      �?             8@52,S
43�       �                 `f�D@����X�?             5@,female�       �                     �?��
ц��?	             *@er (Ali�       �                   �<@�q�q�?             "@ ,"Kalli������������������������       �                      @ 5,,S
43�       �                 `fF<@և���X�?             @ E44,S
4������������������������       �                      @ 20,B96 �       �                 �|Y=@z�G�z�?             @ male,21������������������������       �                     �?(Emily ������������������������       �                     @Mr. Mar������������������������       �                     @ Mr. Jo������������������������       �                      @1,1,2,"������������������������       �                     @1,F.C.C�       �                 h"_@      �?             @5769,9.������������������������       �                     @76,7.77������������������������       �                     �?30434,13�       �                    �?V������?            �B@ ,65306,�       �                    �?�<ݚ�?             "@33638,8�       �                    ;@      �?              @female,�       �                    �?���Q��?             @r",male�       �                 8�T@      �?             @ herine"������������������������       �                      @thur Go������������������������       �                      @ Edwy Ar������������������������       �                     �?r. Ingv������������������������       �                     @an, Mr.������������������������       �                     �? 1,1,"Go�       �                    )@��X��?             <@ 55,0,3,������������������������       �                     @ "Jalsev�       �                 `fFJ@�����?             5@t, Mr. ������������������������       �        
             .@nyon, Mr�       �                     �?�q�q�?             @459,1,2�       �                    7@�q�q�?             @ 
460,0,������������������������       �                     �? 1,"Ande������������������������       �                      @ orley, ������������������������       �                     @ Arthur������������������������       �                     8@ acob Ch�       �                     �?z�G�z�?             @imon",m������������������������       �                     @ Estansl������������������������       �                     �?bell, Mr�                          �?�?�P�a�?(             N@ Montgo�       �                    H@r�q��?             E@ames",m�       �                    �?`2U0*��?             9@rbara",�       �                    �?      �?	             0@ r",male������������������������       �                     �?0,31508�       �                   �F@��S�ۿ?             .@ th)",fe�       �                 `fF:@r�q��?             @ n S (Ma������������������������       �                     @ 917,D,C������������������������       ��q�q�?             @,9.8375������������������������       �                     "@5,52,A1������������������������       �                     "@ 1,,S
47�                       �5L@ҳ�wY;�?             1@,,S
479�                        i?@������?
             .@8,,S
48�       �                 `fF:@���|���?             &@ 2875,,S������������������������       �                     @144,46.�       �                    �?      �?              @ ,0,2398������������������������       �                     �? 5 3594,                          L@և���X�?             @ 34,9.58������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     2@        �t�bh�h*h-K ��h/��R�(KMKK��h]�BP       �{@     �p@     �K@     �h@     �E@      h@     �D@     �g@      @@     �\@              ,@      @@     @Y@      @              :@     @Y@      �?      I@              4@      �?      >@      �?      3@      �?      @      �?      �?              �?      �?                       @              0@              &@      9@     �I@      1@     �G@       @      A@              4@       @      ,@      @      �?              �?      @              @      *@               @      @      &@      @      &@      @       @               @      @                      "@       @              "@      *@      @      "@               @      @      @      @      @      @       @      �?       @      �?                       @       @                      @              �?      @      @      @      �?      @      �?       @              �?      �?              �?      �?              @                      @       @      @      @      �?      @      �?      @                      �?      �?              @      @               @      @      �?       @               @      �?              �?       @              "@      S@       @      H@              ;@       @      5@       @       @      �?      @      �?                      @      @       @      @       @      @       @      @                       @      �?              @                      *@      �?      <@              7@      �?      @              @      �?               @      �?       @                      �?      (@      @              @      (@      �?      (@                      �?     @x@     �Q@     `p@      =@      F@      ,@              "@      F@      @      "@      @      @      @      @                      @      @             �A@       @      .@              4@       @      @              0@       @      "@       @      @       @      @              @             @k@      .@     `j@      *@     �d@      @      N@      �?      $@              I@      �?      0@      �?      0@                      �?      A@             �Z@      @     @Y@      @      3@      @      &@               @      @      @               @      @      �?      @               @      �?      �?      �?             �T@      @     �B@             �F@      @      @@      @      :@       @      7@       @       @       @      5@              @              @      �?              �?      @              *@              @             �F@      @      A@      @      A@      @      5@      �?      @      �?       @               @      �?      1@              *@      @      "@      @      @              @      @               @      @       @      @               @       @               @       @              @                      �?      &@              @       @       @              @       @      @       @               @      @               @             �_@      E@     @R@     �A@      R@      ?@              @      R@      :@      H@      :@      6@      .@      5@      (@      @      @      @       @      �?       @      �?                       @      @              �?      �?      �?                      �?      .@      "@      .@      @      @      @      @      @               @      @      @       @              �?      @      �?                      @      @               @                      @      �?      @              @      �?              :@      &@      @       @      @       @      @       @       @       @               @       @              �?              @              �?              3@      "@              @      3@       @      .@              @       @      �?       @      �?                       @      @              8@              �?      @              @      �?             �J@      @     �A@      @      8@      �?      .@      �?      �?              ,@      �?      @      �?      @               @      �?      "@              "@              &@      @      &@      @      @      @      @              @      @      �?              @      @              @      @              @                       @      2@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ���EhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�G         r                     @�����?�           8�@                                   �?yÏP�?�            �t@ 41m=[3                        03�<@@+K&:~�?[             c@ �P�X                             �?Xny��?(            �N@�P�X                            �H@>A�F<�?             C@                                  �?�t����?             A@                                 @B@�nkK�?             7@       ������������������������       �                     2@        	       
                   �,@z�G�z�?             @ (Y�X  ������������������������       �                     �?"Y�X  ������������������������       �                     @�2Y�X                             �?���!pc�?             &@ +Y�X  ������������������������       �                     �?�2Y�X                            �;@�z�G��?             $@ 0Y�X                            �7@�q�q�?             @        ������������������������       �                      @0$Y�X  ������������������������       �                     �?�X                             D@؇���X�?             @��X  ������������������������       �                     @P��X  ������������������������       �                     �?��X                             �?      �?             @ ��X  ������������������������       �                      @ ��X                            �J@      �?              @ ��X  ������������������������       �                     �?��X  ������������������������       �                     �?��X  ������������������������       �                     7@ ��X  ������������������������       �        3            �V@P��X         =                    �?:���١�?p             f@ ��X         8                     �?�[�IJ�?            �G@��X         5                    �?      �?             C@��X                           ��";@��>4և�?             <@ ��X  ������������������������       �                      @ ��X  !       4                 �̾w@$��m��?             :@     @"       '                 �|Y<@`�Q��?             9@      @#       &                    �?      �?              @       $       %                  �}S@և���X�?             @     @������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?      @(       3                    �?@�0�!��?             1@       )       2                 p�i@@�θ�?	             *@     @*       /                   �A@և���X�?             @      @+       ,                 ���<@      �?             @        ������������������������       �                      @       @-       .                 ��2>@      �?              @       @������������������������       �                     �?     �A@������������������������       �                     �?      :@0       1                  �>@�q�q�?             @       @������������������������       �                     �?        ������������������������       �                      @      "@������������������������       �                     @       @������������������������       �                     @        ������������������������       �                     �?      @6       7                 ��>Y@z�G�z�?             $@     &@������������������������       �                      @       @������������������������       �                      @        9       :                    �?�����H�?             "@      @������������������������       �                     @        ;       <                 pV�C@      �?              @      @������������������������       �                     �?      @������������������������       �                     �?      �?>       m                    �?
�e4���?Q             `@       ?       Z                     �?d�X^_�?I            �\@      @@       O                    B@H.�!���?!             I@      @A       N                 `f�D@�LQ�1	�?             7@      @B       C                 ��I*@��S���?
             .@        ������������������������       �                     @        D       E                   �<@z�G�z�?             $@        ������������������������       �                     @        F       M                   @>@����X�?             @       G       L                 �|�?@���Q��?             @       H       I                 �|Y=@�q�q�?             @        ������������������������       �                     �?        J       K                 `fF<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        P       Y                 ���[@�����H�?             ;@       Q       X                    �?$�q-�?             :@       R       W                 `f�;@�C��2(�?             6@       S       V                   �K@r�q��?             (@        T       U                 ��:@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                     �?        [       l                    �?P�2E��?(            @P@       \       k                   �*@�X�<ݺ?              K@       ]       ^                   �(@$�q-�?            �C@        ������������������������       �        	             ,@        _       `                 �|�<@H%u��?             9@        ������������������������       �                     "@        a       b                 �|�=@     ��?             0@        ������������������������       �                     �?        c       j                   �F@�r����?
             .@       d       i                   @D@z�G�z�?             $@       e       f                    @@�����H�?             "@        ������������������������       �                     @        g       h                   �A@r�q��?             @        ������������������������       ��q�q�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        ������������������������       �                     &@        n       o                    :@X�Cc�?             ,@        ������������������������       �                     @        p       q                    5@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        s                          @l���`��?�            �w@       t       �                    �?B�>�;Q�?�            �w@       u       �                    �?C؇eY�?�            �p@        v                        P��@�ucQ?-�?3            @U@        w       ~                 ���@      �?             8@       x       y                 03S@z�G�z�?
             .@        ������������������������       �                     �?        z       {                   �7@d}h���?	             ,@        ������������������������       �                      @        |       }                    �?�8��8��?             (@        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     "@        �       �                    �?��7��?#            �N@       �       �                 �|Y=@\X��t�?             G@        �       �                    �?     ��?	             0@        �       �                   �2@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?r�q��?             (@       ������������������������       �                      @        �       �                    ;@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?�������?             >@        ������������������������       �                     @        �       �                 @a'@8����?             7@       �       �                 `�j@�q�q�?             5@       �       �                 X��A@�z�G��?             4@       �       �                 �;@�����?             3@       �       �                 03@�q�q�?             2@       �       �                 ��@�t����?             1@        �       �                    �?      �?              @        ������������������������       �                     �?       ������������������������       �                     �?        �       �                 ���@������?	             .@        ������������������������       �                     �?        �       �                    �?����X�?             ,@        ������������������������       �                     @       ������������������������       �                     $@        ������������������������       �                     �?       ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?       ������������������������       �                      @        �       �                    �?z�G�z�?             .@        �       �                    &@      �?              @        ������������������������       �                      @       ������������������������       �                     @       �       �                 ���&@؇���X�?             @        ������������������������       �                     @        �       �                 �|Y=@      �?             @        ������������������������       �                     �?       ������������������������       �                     @        �       �                   �0@X��Oԣ�?t            @g@        ������������������������       �                     @       �       �                    �?�8��8��?o            �f@        �       �                 ���@�q�q�?
             .@        ������������������������       �                     �?        �       �                 �|�;@����X�?	             ,@       �       �                   �9@���|���?             &@       �       �                    8@�<ݚ�?             "@       �       �                   �6@����X�?             @       �       �                  �#@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @       ������������������������       �                      @        ������������������������       �                     @       �       �                 �?�@�FVQ&�?e            �d@        �       �                 �|Y=@`<)�+�?1            @S@       �       �                   �8@p���?             I@       �       �                   �7@ ��WV�?             :@       ������������������������       �                     7@        �       �                 `fF@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     8@        �       �                 �|Y>@�>����?             ;@        �       �                  sW@�t����?
             1@        �       �                 ��,@�q�q�?             @        ������������������������       �                     @        ������������������������       ��q�q�?             @       ������������������������       �                     &@        ������������������������       �        
             $@       �       �                   �3@`���i��?4             V@        �       �                   �1@�θ�?             *@        ������������������������       �                      @       �       �                 `�8"@���!pc�?             &@       �       �                   �2@և���X�?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @       ������������������������       �                     @        �       �                   �:@Х-��ٹ?-            �R@        ������������������������       �                     <@        �       �                   �;@dP-���?             �G@        ������������������������       �                     �?        �       �                 @3�@���.�6�?             G@        �       �                   �?@�q�q�?             @        ������������������������       �                     �?       ������������������������       �                      @        �       �                 ��) @ �#�Ѵ�?            �E@        ������������������������       �                     7@        �       �                 �|�>@ףp=
�?             4@       �       �                 pf� @r�q��?
             (@        ������������������������       �                     �?        �       �                    (@�C��2(�?	             &@        �       �                 �|Y=@z�G�z�?             @        �       �                 ���"@      �?              @        ������������������������       �                     �?       ������������������������       �                     �?       ������������������������       �                     @       ������������������������       �                     @       ������������������������       �                      @       �                          �?������?L             [@       �       �                    �?�BE����?)             O@        �       �                    �?      �?             $@       �       �                    �?X�<ݚ�?             "@       �       �                  S�-@����X�?             @        �       �                 03�)@�q�q�?             @        ������������������������       �                     �?       ������������������������       �                      @       ������������������������       �                     @       ������������������������       �                      @       ������������������������       �                     �?       �       �                    �?�	j*D�?!             J@       �       �                   �3@�P�*�?             ?@        ������������������������       �                     @        �       �                 �|Y=@�q�q�?             ;@        ������������������������       �                     *@       �       �                 03�1@X�Cc�?             ,@        �       �                 ���.@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        �                          �?؇���X�?             5@       �                          �?�KM�]�?             3@       �                        ��y'@�8��8��?	             (@        �       �                 P�@z�G�z�?             @       ������������������������       �                     @       ������������������������       �                     �?        ������������������������       �                     @                                 $@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                                 +@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?*
;&���?#             G@        	                      ��*4@��<b���?             7@        
                        �1@      �?             @        ������������������������       �                      @                                 @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 @�KM�]�?             3@                                 @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@                                 �?���}<S�?             7@       ������������������������       �                     *@                                 @z�G�z�?             $@                              pf�C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                 �?      �?             @        ������������������������       �                     �?                              pf�C@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h*h-K ��h/��R�(KMKK��h]�B�       �{@     �p@     �a@     �g@      @      b@      @      K@      @      ?@      @      >@      �?      6@              2@      �?      @      �?                      @      @       @              �?      @      @       @      �?       @                      �?      �?      @              @      �?              @      �?       @              �?      �?              �?      �?                      7@             �V@     �`@     �E@      ;@      4@      3@      3@      1@      &@               @      1@      "@      1@       @      @      @      @      @              @      @                      �?      ,@      @      $@      @      @      @      @      �?       @              �?      �?              �?      �?              �?       @      �?                       @      @              @                      �?       @       @               @       @               @      �?      @              �?      �?              �?      �?             �Z@      7@     @Y@      ,@     �C@      &@      .@       @      @       @      @               @       @              @       @      @       @      @       @      �?      �?              �?      �?      �?                      �?               @               @       @              8@      @      8@       @      4@       @      $@       @      @       @      @                       @      @              $@              @                      �?      O@      @     �I@      @      B@      @      ,@              6@      @      "@              *@      @              �?      *@       @       @       @       @      �?      @              @      �?       @      �?      @                      �?      @              .@              &@              @      "@              @      @       @               @      @              s@     @S@      s@     �R@      l@     �G@     �M@      :@      5@      @      (@      @      �?              &@      @               @      &@      �?              �?      &@              "@              C@      7@      :@      4@      @      *@      �?      @      �?                      @       @      $@               @       @       @       @                       @      7@      @      @              0@      @      ,@      @      ,@      @      *@      @      (@      @      (@      @      �?      �?              �?      �?              &@      @      �?              $@      @              @      $@                      �?      �?              �?                      �?       @              (@      @      @       @               @      @              @      �?      @              @      �?              �?      @             �d@      5@              @     �d@      .@      $@      @              �?      $@      @      @      @      @       @      @       @      @      �?      @                      �?              �?       @                       @      @             `c@      $@     �R@      @     �H@      �?      9@      �?      7@               @      �?              �?       @              8@              9@       @      .@       @      @       @      @              �?       @      &@              $@             @T@      @      $@      @       @               @      @      @      @              �?      @       @      @             �Q@      @      <@             �E@      @              �?     �E@      @       @      �?              �?       @             �D@       @      7@              2@       @      $@       @              �?      $@      �?      @      �?      �?      �?      �?                      �?      @              @               @              T@      <@     �D@      5@      @      @      @      @       @      @       @      �?              �?       @                      @       @              �?              B@      0@      2@      *@              @      2@      "@      *@              @      "@      �?      "@      �?                      "@      @              2@      @      1@       @      &@      �?      @      �?      @                      �?      @              @      �?              �?      @              �?      �?              �?      �?             �C@      @      2@      @      �?      @               @      �?      �?      �?                      �?      1@       @      �?       @      �?                       @      0@              5@       @      *@               @       @      �?       @               @      �?              @               @       @      �?              �?       @               @      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ:9)bhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMhuh*h-K ��h/��R�(KM��h|�B�G         �                     @e�L��?�           8�@               Y                     �?x@����?�            �u@  l            P                   �J@���(�_�?k            �e@     @                        `V�9@�ӭ�a�?Y             b@     @j@������������������������       �                     @                                  �7@�:���?T             a@        ������������������������       �                     3@               %                   �?@�k��(A�?I            �]@        	                         x;K@Fx$(�?             I@       
                          �<@|��?���?             ;@        ������������������������       �                      @                                  �>@�����?             3@                               �|Y=@���Q��?	             .@        ������������������������       �                      @                                  �<@��
ц��?             *@        ������������������������       �                     @                                  @D@���Q��?             $@ �X  ������������������������       �                     @��X                            �I@z�G�z�?             @ ��X  ������������������������       �                      @��X                             �?�q�q�?             @ ��X  ������������������������       �                      @ ��X  ������������������������       �                     �? ��X  ������������������������       �                     @��X         "                    �?��+7��?             7@��X                             �?�t����?             1@��X  ������������������������       �                     (@P��X                          `f�N@���Q��?             @ ��X  ������������������������       �                      @��X         !                    �?�q�q�?             @��X                            �}S@      �?              @ ��X  ������������������������       �                     �? ��X  ������������������������       �                     �?        ������������������������       �                     �?       @#       $                    �?�q�q�?             @       ������������������������       �                     @      @������������������������       �                      @      �?&       E                 x5Q@�M���?*             Q@     @'       D                 0��M@ҳ�wY;�?             A@       (       1                 ���;@¦	^_�?             ?@      @)       *                 03k:@8�Z$���?             *@      �?������������������������       �                     @        +       ,                    �?z�G�z�?             $@      @������������������������       �                     �?       @-       .                   �C@�<ݚ�?             "@      �?������������������������       �                     @        /       0                    H@�q�q�?             @     �?������������������������       �      �?             @        ������������������������       �                      @       @2       5                    �?b�2�tk�?             2@        3       4                 ��A@      �?              @      @������������������������       �                      @        ������������������������       �                     @      �?6       ;                    �?      �?             $@        7       :                    �?      �?             @      @8       9                    C@�q�q�?             @      �?������������������������       �                      @        ������������������������       �                     �?      @������������������������       �                     �?      �?<       =                   �C@      �?             @        ������������������������       �                     �?      "@>       A                    �?���Q��?             @        ?       @                   @A@      �?              @       @������������������������       �                     �?      �?������������������������       �                     �?        B       C                 �K@�q�q�?             @      @������������������������       �                      @      �?������������������������       �                     �?       @������������������������       �                     @       @F       G                    �?l��\��?             A@      @������������������������       �        
             0@        H       I                    �?r�q��?	             2@        ������������������������       �                      @        J       O                    �?�z�G��?             $@       K       N                 Ј�U@      �?              @        L       M                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        Q       R                 �U'Q@ܷ��?��?             =@       ������������������������       �                     6@        S       T                    �?և���X�?             @        ������������������������       �                      @        U       V                   �K@z�G�z�?             @        ������������������������       �                      @        W       X                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        Z       _                   �1@և���X�?k            �e@        [       \                    �?�}�+r��?             3@       ������������������������       �                     ,@        ]       ^                    #@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        `       �                    L@����3��?_            �c@       a       |                    �?Fx$(�?Y            �b@        b       {                    :@��ϭ�*�?'             M@       c       d                    �?�����H�?            �F@        ������������������������       �                     @        e       z                    �?,���i�?            �D@       f       s                    �?6YE�t�?            �@@       g       j                   �9@�C��2(�?             6@        h       i                   �3@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        k       l                   �'@�}�+r��?             3@        ������������������������       �                     @        m       r                   �,@�8��8��?             (@       n       o                    B@�����H�?             "@       ������������������������       �                     @        p       q                    D@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        t       y                   �E@���!pc�?             &@       u       x                   �;@�����H�?             "@        v       w                   �7@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             *@        }       ~                 �|Y=@�nkK�?2             W@        ������������������������       �                     A@               �                   �*@ 	��p�?!             M@       �       �                    �?(N:!���?            �A@        ������������������������       �                     @,male,32�       �                 �|�=@      �?             @@ male,32�       �                    @�q�q�?             "@nd",mal������������������������       �                     @ter. Eli������������������������       �                     @rtin",ma�       �                   @D@�nkK�?             7@",male,������������������������       �                     &@ale,,1,1�       �                 `f�)@�8��8��?             (@ 5,0,0,3������������������������       �                      @0,349241�       �                   �F@ףp=
�?             $@ 20,0,0,������������������������       ��q�q�?             @er A (Gr������������������������       �                     @1,2,"Wei������������������������       �                     7@0,228414������������������������       �                     @0,0,C.A.�       �                    @��,?S�?�            �v@ PARIS 2�       �                    @$��m��?             :@ ale,19,������������������������       �                     &@eath",ma�       �                    @���Q��?             .@",male,������������������������       �                     @24,0,0,P�       �                    �?      �?              @ ",femal������������������������       �                      @",female�       �                 ��T?@�q�q�?             @ ietari ������������������������       �                      @85,,S
14������������������������       �                     @45,0,2,"�       �                    �?�B���?�            u@ 6,0,2,"�       �                   @C@     ��?=             X@5,,S
14�       �                    �?V�K/��?5            �S@ le,27,0�       �                    �?���B���?             :@Ruby"""�       �                    �?P���Q�?             4@  Michel�       �                 ���,@      �?             @0,2,"By������������������������       �                     @S
151,0,������������������������       �                     �?2.525,,S������������������������       �                     0@,0,11377�       �                 `�@1@�q�q�?             @ 11206,�       �                    �?z�G�z�?             @ .5,0,2,������������������������       �                      @,0,Fa 26�       �                 �|Y=@�q�q�?             @ ,51,0,1������������������������       �                     �?"Katie""������������������������       �                      @",male,3������������������������       �                     �?le",male�       �                   @A@Fmq��?             �J@y",male�       �                   @1@���Q �?            �H@",male,�       �                    �?)O���?             B@h ""Bes�       �                   �5@8�A�0��?             6@ 3,0,3,"�       �                   �3@؇���X�?             @64,0,3,�       �                   !@      �?              @ anula, ������������������������       �                     �?1,3,"Gol������������������������       �                     �?,2,36329������������������������       �                     @an)",fem�       �                 �|�=@��S���?             .@na Bern�       �                 ��&@�n_Y�K�?
             *@Baumann�       �                    ;@���!pc�?             &@ Mr. Le�       �                 03�!@և���X�?             @ Wyckof�       �                   �7@      �?             @ rthur",������������������������       �                      @nor Ilee�       �                 pff@      �?              @ tti Wil������������������������       �                     �?ith, Mr.������������������������       �                     �?lasen, M������������������������       �                     @ebre, Ma������������������������       �                     @sham, Mi������������������������       �                      @179,0,2,������������������������       �                      @eonard, �       �                    �?����X�?             ,@nstance�       �                    �?�θ�?             *@r. Rene�       �                 ���)@�q�q�?             "@ er. Cla������������������������       �                     @"Becker,�       �                 �|�;@      �?             @ nk-Heil������������������������       �                     �?S
186,0,������������������������       �                     @1,3,"O'B������������������������       �                     @1,0,3703������������������������       �                     �? Rolmane������������������������       �        	             *@hn",male������������������������       �                     @e,36,0,0������������������������       �                     1@2,0,0,23�                          �?P�_��I�?�             n@424,13,�       �                    �?      �?�             l@ ne",fem�       �                 �=/@�<ݚ�?$             K@chel M"�       �                   �7@@�0�!��?"            �I@ eph (Ma�       �                    �?      �?             @1,"Lure������������������������       �                      @197,0,3,������������������������       �                      @Olsen, M�       �                    �?��0{9�?            �G@ 1,3,"Ma�       �                    �?�X�<ݺ?             2@,,Q
200�       �                 �|Y?@��S�ۿ?             .@,0,0,24�       �                 �|Y;@�����H�?             "@ 28,0,0,������������������������       �                     �?. 2343,6�       �                 ���@      �?              @ 3101264������������������������       �                     @2628,7.2�       �                 p&�@      �?             @5 3540,������������������������       ��q�q�?             @1,347054������������������������       �                     �?32,1,0,3������������������������       �                     @le,26,0,������������������������       �                     @female,1�       �                  ��@V�a�� �?             =@ ,0,1122������������������������       �                     @.Q. 3101�       �                    �?���!pc�?             6@5,0,0,F�       �                 X��A@����X�?             5@2,0,0,A�       �                   @'@ҳ�wY;�?	             1@le,30,0������������������������       �      �?             0@367229,7������������������������       �                     �?5273,113������������������������       �                     @0,STON/O������������������������       �                     �?l",male,������������������������       �                     @le,32,0,�       �                   �0@��O���?q            @e@ 0,0,0,W�       �                 pf�@      �?             @ ,male,1������������������������       �                     �?s H",mal�       �                    �?���Q��?             @ale,51,�       �                 pFD!@      �?             @ 0,34923������������������������       �                      @38,1,0,1������������������������       �                      @e,22,0,0������������������������       �                     �?e,19,0,0�                         @@@���C"��?l            �d@y"")",m�                          �? �	.��?V            ``@ne Jona�                       �!&B@�|K��2�?U             `@lde",fe�                       �|�=@�[|x��?S            �_@khardt �                       �|Y=@@-�_ .�?K            �[@,"Larss�                          �?�F��O�?7            @R@"Sjoste�       �                   �:@�U�=���?1            �P@Asplund�       �                 @3�@@9G��?'            �H@35,0,2,������������������������       �                     :@66,10.5,�       �                 0S5 @���}<S�?             7@ C. 6609�       �                   �2@      �?              @ ,,S
238������������������������       �                     �?.A. 3192�       �                   �3@؇���X�?             @ ,19,0,0������������������������       ��q�q�?             @0,0,SCO/������������������������       �                     @,1,0,266������������������������       �                     .@female,,                       pf� @@�0�!��?
             1@es",mal������������������������       �                     "@                              ���)@      �?              @                               �;@      �?             @        ������������������������       �                      @                                �<@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        	                         5@؇���X�?             @        
                      �Y�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     C@                                �?@������?             .@                                �>@      �?              @                              (Se!@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @                              pff@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                 �?؇���X�?             @                             ��I @r�q��?             @       ������������������������       �      �?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �@@        ������������������������       �        	             1@        �t�b�(z      h�h*h-K ��h/��R�(KMKK��h]�B�       �{@     �p@     �d@     �f@     �P@     �Z@     �D@     �Y@      @              A@     �Y@              3@      A@      U@      3@      ?@      *@      ,@               @      *@      @      "@      @       @              @      @      @              @      @              @      @      �?       @               @      �?       @                      �?      @              @      1@       @      .@              (@       @      @               @       @      �?      �?      �?              �?      �?              �?              @       @      @                       @      .@     �J@      (@      6@      "@      6@       @      &@              @       @       @              �?       @      @              @       @      @       @       @               @      @      &@       @      @       @                      @      @      @       @       @       @      �?       @                      �?              �?      @      @      �?               @      @      �?      �?              �?      �?              �?       @               @      �?              @              @      ?@              0@      @      .@               @      @      @      �?      @      �?      @              @      �?                      @       @              :@      @      6@              @      @               @      @      �?       @               @      �?              �?       @              Y@     �R@      �?      2@              ,@      �?      @              @      �?             �X@     �L@     @W@     �L@      @     �J@      @      D@              @      @      B@      @      <@       @      4@      �?       @      �?                       @      �?      2@              @      �?      &@      �?       @              @      �?       @      �?                       @              @      @       @      �?       @      �?      @      �?                      @              @       @                       @              *@      V@      @      A@              K@      @      ?@      @      @              <@      @      @      @      @                      @      6@      �?      &@              &@      �?       @              "@      �?       @      �?      @              7@              @             @q@     �U@      "@      1@              &@      "@      @      @               @      @               @       @      @       @                      @     �p@     �Q@      K@      E@     �B@      E@      @      5@      �?      3@      �?      @              @      �?                      0@      @       @      @      �?       @               @      �?              �?       @                      �?      @@      5@      @@      1@      3@      1@      "@      *@      �?      @      �?      �?      �?                      �?              @       @      @       @      @       @      @      @      @      �?      @               @      �?      �?      �?                      �?      @              @                       @               @      $@      @      $@      @      @      @      @              �?      @      �?                      @      @                      �?      *@                      @      1@             �j@      <@     �h@      <@      E@      (@      E@      "@       @       @               @       @              D@      @      1@      �?      ,@      �?       @      �?      �?              @      �?      @              @      �?       @      �?      �?              @              @              7@      @      @              0@      @      .@      @      &@      @      $@      @      �?              @              �?                      @     @c@      0@      @      @      �?               @      @       @       @               @       @                      �?     �b@      *@     �]@      *@      ]@      *@      ]@      $@     @Z@      @     �P@      @     �N@      @     �G@       @      :@              5@       @      @       @              �?      @      �?       @      �?      @              .@              ,@      @      "@              @      @      �?      @               @      �?      �?      �?                      �?      @              @      �?      �?      �?      �?                      �?      @              C@              &@      @      @      @      @       @      @                       @       @      �?       @                      �?      @      �?      @      �?      @      �?       @              �?                      @       @             �@@              1@        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh&hNhJ�BHzhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtMIhuh*h-K ��h/��R�(KMI��h|�B@R         N                    �?�t����?�           8�@                                   �?�9��L~�?^            �b@                                `�@1@�C��2(�?)            �P@      @                           �?�E��ӭ�?             2@                                  �?�8��8��?             (@       ������������������������       �                     @                                P��+@z�G�z�?             @        ������������������������       �                      @        	       
                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?�q�q�?             @     @                        �&�)@���Q��?             @      @������������������������       �                     �?      �?                          �-@      �?             @        ������������������������       �                      @      �?                        ���,@      �?              @      @������������������������       �                     �?      .@������������������������       �                     �?      (@������������������������       �                     �?      �?                          �H@@��8��?             H@     @������������������������       �                     D@                                   �?      �?              @                                   �?      �?             @                               ,w�U@�q�q�?             @      @������������������������       �                     �?        ������������������������       �                      @      �?������������������������       �                     �?      @������������������������       �                     @     �D@       -                 pF�#@�t����?5            @U@      @       "                   �5@�#-���?            �A@                !                 �{@      �?              @       @������������������������       �                     �?        ������������������������       �                     �?      �?#       $                 ���@�FVQ&�?            �@@        ������������������������       �                     ,@      1@%       (                 �|Y=@�KM�]�?             3@      @&       '                   @@      �?             @     @������������������������       �                     @      5@������������������������       �                     �?        )       ,                   @@��S�ۿ?
             .@        *       +                 �|�=@z�G�z�?             @     �?������������������������       �      �?             @      *@������������������������       �                     �?      �?������������������������       �                     $@      @.       I                     @� �	��?             I@     �?/       D                     �?�D����?             E@       0       C                   �H@X�<ݚ�?             B@     @1       2                 �|Y<@���!pc�?             6@        ������������������������       �                     @        3       >                    �?ҳ�wY;�?             1@     <@4       ;                 `f�A@�q�q�?             (@      @5       :                 X�,@@      �?              @     �?6       7                 �ܵ<@���Q��?             @        ������������������������       �                     �?        8       9                 ��2>@      �?             @      @������������������������       �                     @        ������������������������       �                     �?      0@������������������������       �                     @       @<       =                 @�Cq@      �?             @     *@������������������������       �                     @      @������������������������       �                     �?        ?       @                   @H@z�G�z�?             @      �?������������������������       �                     �?      @A       B                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ,@        E       F                 ���@@r�q��?             @       ������������������������       �                     @        G       H                    �?      �?              @        ������������������������       �                     �?       ������������������������       �                     �?       J       M                    �?      �?              @        K       L                   �3@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        O       �                   �3@�钹H��?^           ��@        P       �                    @��o	��?D             ]@       Q       v                    �?8�$�>�?4            �U@       R       S                    �?
;&����?             G@        ������������������������       �                     @        T       q                    6@�G��l��?             E@       U       n                    �?���Q��?            �A@       V       ]                    �?J�8���?             =@        W       X                   �1@z�G�z�?             @        ������������������������       �                     �?       Y       \                 ��!@      �?             @       Z       [                 P��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @       ^       a                     @      �?             8@        _       `                   �2@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        b       g                   �1@���y4F�?             3@        c       f                   �0@      �?              @        d       e                 pf�@�q�q�?             @        ������������������������       �                     �?       ������������������������       �      �?              @        ������������������������       �                     @        h       m                 0S5 @���!pc�?             &@        i       j                   �2@      �?             @        ������������������������       �                      @       k       l                 �?�@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        o       p                   �2@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        r       s                     �?؇���X�?             @        ������������������������       �                     �?       t       u                   �1@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        w       ~                    �?z�G�z�?             D@        x       y                     @�t����?             1@       ������������������������       �                     $@       z       {                    �?����X�?             @        ������������������������       �                     @        |       }                 `f7@      �?             @       ������������������������       �                      @        ������������������������       �                      @              �                    )@��+7��?             7@       �       �                    �?�KM�]�?             3@       ������������������������       �                     *@        �       �                    �?�q�q�?             @       �       �                    �?z�G�z�?             @        ������������������������       �                     @        �       �                     �?      �?              @        ������������������������       �                     �?       ������������������������       �                     �?       ������������������������       �                     �?       ������������������������       �                     @        �       �                    �?z�G�z�?             >@        �       �                    @ҳ�wY;�?             1@        ������������������������       �                     @        �       �                    *@��
ц��?             *@       �       �                    @�z�G��?             $@        �       �                    @      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             *@        �       �                     @�/e�U��?           �{@        �       �                    �?      �?v             g@       �       �                    �?*��w\��?\            �b@        �       �                    :@=QcG��?            �G@        �       �                   �3@���Q��?             @        ������������������������       �                      @       ������������������������       �                     @        �       �                   �B@�Ń��̧?             E@       ������������������������       �                     9@        �       �                   @C@�IєX�?             1@        ������������������������       �                     �?        ������������������������       �        
             0@        �       �                    �?��[�8��?B            �Y@        ������������������������       �                     �?       �       �                     �?�C+����?A            @Y@       �       �                    �?���Q �?!            �H@       �       �                   �B@�z�G��?             D@       �       �                   �A@���Q��?             >@       �       �                   �>@�q�q�?             ;@       �       �                   @>@և���X�?             5@       �       �                 �̌*@�q�q�?             2@        ������������������������       �                     @        �       �                 `fF<@և���X�?
             ,@       �       �                   @L@�eP*L��?             &@       �       �                    H@      �?              @       �       �                 �|�<@      �?             @        ������������������������       �                     �?        �       �                 �|�?@���Q��?             @        ������������������������       �                     �?       �       �                   �C@      �?             @        ������������������������       �                     �?        ������������������������       ��q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        �       �                 �|Y=@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        �       �                    =@X�<ݚ�?             "@        ������������������������       �                     �?        �       �                 ��<R@      �?              @       �       �                   �C@z�G�z�?             @        ������������������������       �                      @        �       �                  x#J@�q�q�?             @        ������������������������       �                     �?        �       �                 �K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    ,@4��?�?              J@       �       �                 `f�)@�חF�P�?             ?@        ������������������������       �        	             (@        �       �                   �A@�d�����?             3@        �       �                 �|Y<@      �?              @        ������������������������       �                      @        �       �                 �|�=@�q�q�?             @        ������������������������       �                     �?        �       �                    @@���Q��?             @        ������������������������       �                     �?       ������������������������       �      �?             @        �       �                   �F@�C��2(�?             &@       �       �                   @D@z�G�z�?             @        ������������������������       �                      @        ������������������������       ��q�q�?             @       ������������������������       �                     @        ������������������������       �                     5@        �       �                   �M@��R[s�?            �A@       �       �                    F@     ��?             @@       �       �                    B@�+e�X�?             9@       �       �                    �?R���Q�?             4@       ������������������������       �                     1@       ������������������������       �                     @        �       �                    �?���Q��?             @        ������������������������       �                      @       ������������������������       �                     @       ������������������������       �                     @        ������������������������       �                     @        �                          �?�����D�?�            @p@        �                          �?�ʻ����?.             Q@       �       �                 ��@�~8�e�?$            �I@        �       �                    �?@�0�!��?             1@       �       �                 ���@ףp=
�?             $@        ������������������������       �                     �?       ������������������������       �                     "@       �       �                 pff@����X�?             @       �       �                 �|�9@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�ʻ����?             A@        ������������������������       �                     @       �                         �>@d��0u��?             >@       �       �                 ��&@l��
I��?             ;@       �       �                   �@�r����?
             .@        �       �                 �&B@      �?             @       �       �                   �7@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        �                          4@      �?             (@       �       �                   �:@      �?              @        ������������������������       �                     �?        �                           �?؇���X�?             @        ������������������������       �                     @                                �.@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                              �|�:@�IєX�?
             1@        ������������������������       �                     �?        ������������������������       �        	             0@        	      D                ���5@     ��?v             h@       
      ?                   �?�L���?r             g@             6                ���"@d#,����?e            �d@                                �?@�+9\J�?Z            �b@                              �|Y=@؇���X�?             5@                               ��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                              X�I@�KM�]�?             3@                             ���@�t����?             1@        ������������������������       �                      @                              ��(@�<ݚ�?             "@       ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                      @                                �7@����?K            @`@        ������������������������       �                    �A@                              ���@<����?7            �W@        ������������������������       �        	             2@                                @8@�s�c���?.            @S@                              03@      �?             @        ������������������������       �                      @        ������������������������       �                      @               1                @3�@�F��O�?,            @R@       !      "                �|Y=@X�EQ]N�?            �E@        ������������������������       �                     .@        #      0                  �C@�>4և��?             <@       $      %                pf�@�E��ӭ�?             2@        ������������������������       �                     @        &      /                   B@�q�q�?
             (@       '      .                  @@@���|���?	             &@       (      )                  �@���Q��?             $@        ������������������������       �                     @        *      +                �|�>@؇���X�?             @        ������������������������       �                     @        ,      -                �?�@�q�q�?             @        ������������������������       �                     �?        ������������������������       �      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     $@        2      5                �|Y<@(;L]n�?             >@        3      4                  �:@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ;@        7      <                �|�=@d}h���?             ,@       8      9                  �<@�C��2(�?	             &@       ������������������������       �                     @        :      ;                �|Y=@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        =      >                  �A@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        @      C                pf� @P���Q�?             4@        A      B                ��Y@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             (@        E      H                   �?և���X�?             @        F      G                   �?���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h*h-K ��h/��R�(KMIKK��h]�B�       �z@     �q@     �P@     @U@      @      N@      @      *@      �?      &@              @      �?      @               @      �?       @      �?                       @      @       @      @       @              �?      @      �?       @              �?      �?              �?      �?              �?              �?     �G@              D@      �?      @      �?      @      �?       @      �?                       @              �?              @      N@      9@      @@      @      �?      �?      �?                      �?      ?@       @      ,@              1@       @      @      �?      @                      �?      ,@      �?      @      �?      @      �?      �?              $@              <@      6@      9@      1@      4@      0@      @      0@              @      @      &@      @      @       @      @       @      @      �?              �?      @              @      �?                      @      @      �?      @                      �?      �?      @              �?      �?      @              @      �?              ,@              @      �?      @              �?      �?              �?      �?              @      @      @       @               @      @                      @     `v@     @i@      K@      O@      >@      L@      6@      8@              @      6@      4@      5@      ,@      3@      $@      �?      @              �?      �?      @      �?      �?              �?      �?                       @      2@      @      @       @      @                       @      .@      @      @      �?       @      �?      �?              �?      �?      @               @      @      �?      @               @      �?      �?      �?                      �?      @               @      @       @                      @      �?      @              �?      �?      @      �?                      @       @      @@       @      .@              $@       @      @              @       @       @               @       @              @      1@       @      1@              *@       @      @      �?      @              @      �?      �?      �?                      �?      �?              @              8@      @      &@      @      @              @      @      @      @      �?      @      �?                      @      @                      @      *@              s@     �a@      W@      W@     �T@     �P@      @      F@       @      @       @                      @      �?     �D@              9@      �?      0@      �?                      0@      T@      6@      �?             �S@      6@      @@      1@      <@      (@      2@      (@      2@      "@      (@      "@      (@      @      @               @      @      @      @      @      @      @      @              �?      @       @      �?               @       @              �?       @      �?               @      @               @      �?       @                      �?              @      @                      @      $@              @      @              �?      @      @      @      �?       @               @      �?      �?              �?      �?              �?      �?                      @     �G@      @      :@      @      (@              ,@      @      @      @       @               @      @              �?       @      @      �?              �?      @      $@      �?      @      �?       @               @      �?      @              5@              "@      :@      @      :@      @      3@      @      1@              1@      @              @       @               @      @                      @      @             �j@      H@      C@      >@      6@      =@      @      ,@      �?      "@      �?                      "@       @      @       @       @               @       @                      @      3@      .@              @      3@      &@      3@       @      *@       @       @       @       @      �?              �?       @                      �?      &@              @      @       @      @      �?              �?      @              @      �?      @      �?                      @      @                      @      0@      �?              �?      0@             �e@      2@     @e@      .@     �b@      ,@     �a@      &@      2@      @      �?      �?      �?                      �?      1@       @      .@       @       @              @       @      @       @      �?               @             �^@       @     �A@             �U@       @      2@             @Q@       @       @       @               @       @             �P@      @      C@      @      .@              7@      @      *@      @      @              @      @      @      @      @      @              @      @      �?      @               @      �?      �?              �?      �?      �?                      �?      $@              =@      �?       @      �?       @                      �?      ;@              &@      @      $@      �?      @              @      �?              �?      @              �?       @               @      �?              3@      �?      @      �?      @                      �?      (@              @      @       @      @       @                      @       @        �t�bubhhubehhub.